** sch_path: /home/schippes/.xschem/xschem_library/xschem_sky130/xschem_verilog_import/audiodac.sch
**.subckt audiodac VGND VPWR clk_i ds_n_o ds_o fifo_ack_o fifo_empty_o fifo_full_o fifo_rdy_i mode_i
*+ rst_n_i
*+ fifo_i[15],fifo_i[14],fifo_i[13],fifo_i[12],fifo_i[11],fifo_i[10],fifo_i[9],fifo_i[8],fifo_i[7],fifo_i[6],fifo_i[5],fifo_i[4],fifo_i[3],fifo_i[2],fifo_i[1],fifo_i[0] osr_i[1],osr_i[0] volume_i[3],volume_i[2],volume_i[1],volume_i[0]
*.ipin VGND
*.ipin VPWR
*.ipin clk_i
*.opin ds_n_o
*.opin ds_o
*.opin fifo_ack_o
*.opin fifo_empty_o
*.opin fifo_full_o
*.ipin fifo_rdy_i
*.ipin mode_i
*.ipin rst_n_i
*.ipin
*+ fifo_i[15],fifo_i[14],fifo_i[13],fifo_i[12],fifo_i[11],fifo_i[10],fifo_i[9],fifo_i[8],fifo_i[7],fifo_i[6],fifo_i[5],fifo_i[4],fifo_i[3],fifo_i[2],fifo_i[1],fifo_i[0]
*.ipin osr_i[1],osr_i[0]
*.ipin volume_i[3],volume_i[2],volume_i[1],volume_i[0]
XANTENNA_0 _0091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 _0992_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1011_ fifo_dfifo__reg_o9_c_o14_c VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__inv_2
X_1012_ net21 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__clkbuf_1
X_1013_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__clkbuf_4
X_1014_ fifo_dwrite__ptr_o1_c VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1015_ fifo_dwrite__ptr_o0_c VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1016_ fifo_dwrite__ptr_o1_c VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__inv_2
X_1017_ fifo_dwrite__ptr_o0_c VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__clkinv_2
X_1018_ _0784_ _0785_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__or2_2
X_1019_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__inv_2
X_1020_ fifo_dwrite__ptr_o2_c VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__inv_2
X_1021_ fifo_dwrite__ptr_o3_c VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__inv_2
X_1022_ _0788_ _0786_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__o21a_1
X_1023_ fifo_dwrite__ptr_o2_c _0787_ fifo_dwrite__ptr_o3_c _0790_ VGND VGND VPWR VPWR _0791_
+ sky130_fd_sc_hd__a31o_1
X_1024_ _0786_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__clkbuf_2
X_1025_ _0788_ _0792_ fifo_dwrite__ptr_o2_c _0787_ VGND VGND VPWR VPWR _0793_
+ sky130_fd_sc_hd__o22a_1
X_1026_ net21 VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__inv_2
X_1027_ net17 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__inv_2
X_1028_ fifo_dread__ptr_o3_c VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
X_1029_ _0791_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__inv_2
X_1030_ fifo_dread__ptr_o1_c VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
X_1031_ fifo_dwrite__ptr_o1_c fifo_dwrite__ptr_o0_c _0786_ VGND VGND VPWR VPWR _0797_
+ sky130_fd_sc_hd__o21ai_1
X_1032_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__inv_2
X_1033_ fifo_dread__ptr_o0_c VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__inv_2
X_1034_ fifo_dread__ptr_o0_c _0785_ _0799_ fifo_dwrite__ptr_o0_c VGND VGND VPWR VPWR _0800_
+ sky130_fd_sc_hd__a22o_1
X_1035_ fifo_dread__ptr_o2_c VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
X_1036_ fifo_dread__ptr_o2_c fifo_dwrite__ptr_o2_c _0009_ _0788_ VGND VGND VPWR VPWR _0801_
+ sky130_fd_sc_hd__o22a_1
X_1037_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__inv_2
X_1038_ _0786_ _0801_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__or2_1
X_1039_ fifo_dread__ptr_o1_c _0797_ _0787_ _0802_ _0803_ VGND VGND VPWR VPWR _0804_
+ sky130_fd_sc_hd__o221a_1
X_1040_ _0008_ _0798_ _0800_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__o211a_1
X_1041_ _0010_ _0796_ fifo_dread__ptr_o3_c _0791_ _0805_ VGND VGND VPWR VPWR net30
+ sky130_fd_sc_hd__o221a_1
X_1042_ _0795_ fifo_dfifo__rdy__last net30 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or3_2
X_1043_ _0794_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__or2_1
X_1044_ _0793_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__or2_1
X_1045_ _0791_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or2_1
X_1046_ _0782_ _0783_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__or3_4
X_1047_ _0781_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__nand2_2
X_1048_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__clkbuf_2
X_1049_ _0810_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_2
X_1050_ _0794_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__clkbuf_2
X_1051_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__clkbuf_2
X_1052_ _0806_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1053_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__buf_2
X_1054_ _0815_ _0817_ net6 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__or3b_2
X_1055_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkbuf_2
X_1056_ _0779_ _0812_ _0813_ _0819_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o22ai_1
X_1057_ fifo_dfifo__reg_o9_c_o13_c VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__inv_2
X_1058_ _0815_ _0817_ net5 VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or3b_2
X_1059_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__clkbuf_2
X_1060_ _0820_ _0812_ _0813_ _0822_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o22ai_1
X_1061_ fifo_dfifo__reg_o9_c_o12_c VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__inv_2
X_1062_ _0794_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__buf_2
X_1063_ _0824_ _0817_ net4 VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__or3b_4
X_1064_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__clkbuf_2
X_1065_ _0823_ _0812_ _0813_ _0826_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o22ai_1
X_1066_ fifo_dfifo__reg_o9_c_o11_c VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__inv_2
X_1067_ _0816_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__clkbuf_2
X_1068_ _0824_ _0828_ net3 VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__or3b_4
X_1069_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_2
X_1070_ _0827_ _0812_ _0813_ _0830_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__o22ai_1
X_1071_ fifo_dfifo__reg_o9_c_o10_c VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__inv_2
X_1072_ _0824_ _0828_ net2 VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__or3b_2
X_1073_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__buf_2
X_1074_ _0831_ _0812_ _0813_ _0833_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__o22ai_1
X_1075_ fifo_dfifo__reg_o9_c_o9_c VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__inv_2
X_1076_ _0811_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__buf_2
X_1077_ _0810_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__buf_2
X_1078_ _0824_ _0828_ net16 VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__or3b_2
X_1079_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__clkbuf_2
X_1080_ _0834_ _0835_ _0836_ _0838_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__o22ai_1
X_1081_ fifo_dfifo__reg_o9_c_o8_c VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__inv_2
X_1082_ _0824_ _0828_ net15 VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__or3b_2
X_1083_ _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__buf_2
X_1084_ _0839_ _0835_ _0836_ _0841_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__o22ai_1
X_1085_ fifo_dfifo__reg_o9_c_o7_c VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__inv_2
X_1086_ _0794_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__clkbuf_2
X_1087_ _0843_ _0828_ net14 VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or3b_2
X_1088_ _0844_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__clkbuf_2
X_1089_ _0842_ _0835_ _0836_ _0845_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o22ai_1
X_1090_ fifo_dfifo__reg_o9_c_o6_c VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__inv_2
X_1091_ _0806_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__clkbuf_2
X_1092_ _0843_ _0847_ net13 VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__or3b_2
X_1093_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_2
X_1094_ _0846_ _0835_ _0836_ _0849_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o22ai_1
X_1095_ fifo_dfifo__reg_o9_c_o5_c VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__inv_2
X_1096_ _0843_ _0847_ net12 VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__or3b_4
X_1097_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__clkbuf_2
X_1098_ _0850_ _0835_ _0836_ _0852_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o22ai_1
X_1099_ fifo_dfifo__reg_o9_c_o4_c VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__inv_2
X_1100_ _0811_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_2
X_1101_ _0810_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_2
X_1102_ _0843_ _0847_ net11 VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__or3b_2
X_1103_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__clkbuf_2
X_1104_ _0853_ _0854_ _0855_ _0857_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__o22ai_1
X_1105_ fifo_dfifo__reg_o9_c_o3_c VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__inv_2
X_1106_ _0843_ _0847_ net10 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or3b_4
X_1107_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__clkbuf_2
X_1108_ _0858_ _0854_ _0855_ _0860_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__o22ai_1
X_1109_ fifo_dfifo__reg_o9_c_o2_c VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__inv_2
X_1110_ _0814_ _0847_ net9 VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__or3b_4
X_1111_ _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__clkbuf_2
X_1112_ _0861_ _0854_ _0855_ _0863_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o22ai_1
X_1113_ fifo_dfifo__reg_o9_c_o1_c VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__inv_2
X_1114_ _0814_ _0816_ net8 VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__or3b_4
X_1115_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__clkbuf_2
X_1116_ _0864_ _0854_ _0855_ _0866_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o22ai_1
X_1117_ fifo_dfifo__reg_o9_c_o0_c VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__inv_2
X_1118_ _0814_ _0816_ net1 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__or3b_2
X_1119_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__clkbuf_2
X_1120_ _0867_ _0854_ _0855_ _0869_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__o22ai_1
X_1121_ net21 VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__buf_2
X_1122_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1123_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__buf_2
X_1124_ _0792_ _0809_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2_4
X_1125_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__clkbuf_2
X_1126_ net7 VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__clkbuf_2
X_1127_ _0873_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__clkinv_2
X_1128_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__clkbuf_2
X_1129_ _0872_ _0874_ fifo_dfifo__reg_o8_c_o15_c _0875_ _0877_ VGND VGND VPWR VPWR _0434_
+ sky130_fd_sc_hd__a32o_1
X_1130_ net6 VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__clkbuf_2
X_1131_ _0872_ _0874_ fifo_dfifo__reg_o8_c_o14_c _0878_ _0877_ VGND VGND VPWR VPWR _0433_
+ sky130_fd_sc_hd__a32o_1
X_1132_ _0871_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__clkbuf_2
X_1133_ net5 VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__clkbuf_2
X_1134_ _0879_ _0874_ fifo_dfifo__reg_o8_c_o13_c _0880_ _0877_ VGND VGND VPWR VPWR _0432_
+ sky130_fd_sc_hd__a32o_1
X_1135_ net4 VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_2
X_1136_ _0879_ _0874_ fifo_dfifo__reg_o8_c_o12_c _0881_ _0877_ VGND VGND VPWR VPWR _0431_
+ sky130_fd_sc_hd__a32o_1
X_1137_ net3 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__clkbuf_2
X_1138_ _0879_ _0874_ fifo_dfifo__reg_o8_c_o11_c _0882_ _0877_ VGND VGND VPWR VPWR _0430_
+ sky130_fd_sc_hd__a32o_1
X_1139_ _0873_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__clkbuf_2
X_1140_ net2 VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__buf_2
X_1141_ _0876_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__clkbuf_2
X_1142_ _0879_ _0883_ fifo_dfifo__reg_o8_c_o10_c _0884_ _0885_ VGND VGND VPWR VPWR _0429_
+ sky130_fd_sc_hd__a32o_1
X_1143_ net16 VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__buf_2
X_1144_ _0879_ _0883_ fifo_dfifo__reg_o8_c_o9_c _0886_ _0885_ VGND VGND VPWR VPWR _0428_
+ sky130_fd_sc_hd__a32o_1
X_1145_ _0871_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__clkbuf_2
X_1146_ net15 VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__clkbuf_2
X_1147_ _0887_ _0883_ fifo_dfifo__reg_o8_c_o8_c _0888_ _0885_ VGND VGND VPWR VPWR _0427_
+ sky130_fd_sc_hd__a32o_1
X_1148_ net14 VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__clkbuf_2
X_1149_ _0887_ _0883_ fifo_dfifo__reg_o8_c_o7_c _0889_ _0885_ VGND VGND VPWR VPWR _0426_
+ sky130_fd_sc_hd__a32o_1
X_1150_ net13 VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__clkbuf_2
X_1151_ _0887_ _0883_ fifo_dfifo__reg_o8_c_o6_c _0890_ _0885_ VGND VGND VPWR VPWR _0425_
+ sky130_fd_sc_hd__a32o_1
X_1152_ _0873_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__clkbuf_2
X_1153_ net12 VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__buf_2
X_1154_ _0876_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__clkbuf_2
X_1155_ _0887_ _0891_ fifo_dfifo__reg_o8_c_o5_c _0892_ _0893_ VGND VGND VPWR VPWR _0424_
+ sky130_fd_sc_hd__a32o_1
X_1156_ net11 VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__buf_2
X_1157_ _0887_ _0891_ fifo_dfifo__reg_o8_c_o4_c _0894_ _0893_ VGND VGND VPWR VPWR _0423_
+ sky130_fd_sc_hd__a32o_1
X_1158_ _0870_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1159_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__buf_2
X_1160_ net10 VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__buf_2
X_1161_ _0896_ _0891_ fifo_dfifo__reg_o8_c_o3_c _0897_ _0893_ VGND VGND VPWR VPWR _0422_
+ sky130_fd_sc_hd__a32o_1
X_1162_ net9 VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__buf_2
X_1163_ _0896_ _0891_ fifo_dfifo__reg_o8_c_o2_c _0898_ _0893_ VGND VGND VPWR VPWR _0421_
+ sky130_fd_sc_hd__a32o_1
X_1164_ net8 VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__buf_2
X_1165_ _0896_ _0891_ fifo_dfifo__reg_o8_c_o1_c _0899_ _0893_ VGND VGND VPWR VPWR _0420_
+ sky130_fd_sc_hd__a32o_1
X_1166_ net1 VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__clkbuf_2
X_1167_ _0896_ _0873_ fifo_dfifo__reg_o8_c_o0_c _0900_ _0876_ VGND VGND VPWR VPWR _0419_
+ sky130_fd_sc_hd__a32o_1
X_1168_ fifo_dfifo__reg_o7_c_o15_c VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__inv_2
X_1169_ _0796_ _0807_ _0793_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__or3b_2
X_1170_ _0807_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__buf_2
X_1171_ _0798_ _0903_ _0785_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__o22ai_4
X_1172_ _0902_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__or2_4
X_1173_ _0781_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nand2_4
X_1174_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__clkbuf_2
X_1175_ _0814_ _0816_ net7 VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__or3b_2
X_1176_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__clkbuf_2
X_1177_ _0905_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__clkbuf_2
X_1178_ _0901_ _0907_ _0909_ _0910_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__o22ai_1
X_1179_ fifo_dfifo__reg_o7_c_o14_c VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__inv_2
X_1180_ _0911_ _0907_ _0819_ _0910_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o22ai_1
X_1181_ fifo_dfifo__reg_o7_c_o13_c VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__inv_2
X_1182_ _0912_ _0907_ _0822_ _0910_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__o22ai_1
X_1183_ fifo_dfifo__reg_o7_c_o12_c VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__inv_2
X_1184_ _0913_ _0907_ _0826_ _0910_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o22ai_1
X_1185_ fifo_dfifo__reg_o7_c_o11_c VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__inv_2
X_1186_ _0914_ _0907_ _0830_ _0910_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o22ai_1
X_1187_ fifo_dfifo__reg_o7_c_o10_c VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__inv_2
X_1188_ _0906_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__clkbuf_2
X_1189_ _0905_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__clkbuf_2
X_1190_ _0915_ _0916_ _0833_ _0917_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o22ai_1
X_1191_ fifo_dfifo__reg_o7_c_o9_c VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__inv_2
X_1192_ _0918_ _0916_ _0838_ _0917_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__o22ai_1
X_1193_ fifo_dfifo__reg_o7_c_o8_c VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__inv_2
X_1194_ _0919_ _0916_ _0841_ _0917_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__o22ai_1
X_1195_ fifo_dfifo__reg_o7_c_o7_c VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__inv_2
X_1196_ _0920_ _0916_ _0845_ _0917_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o22ai_1
X_1197_ fifo_dfifo__reg_o7_c_o6_c VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__inv_2
X_1198_ _0921_ _0916_ _0849_ _0917_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__o22ai_1
X_1199_ fifo_dfifo__reg_o7_c_o5_c VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__inv_2
X_1200_ _0906_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__clkbuf_2
X_1201_ _0905_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__clkbuf_2
X_1202_ _0922_ _0923_ _0852_ _0924_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o22ai_1
X_1203_ fifo_dfifo__reg_o7_c_o4_c VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__inv_2
X_1204_ _0925_ _0923_ _0857_ _0924_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o22ai_1
X_1205_ fifo_dfifo__reg_o7_c_o3_c VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__inv_2
X_1206_ _0926_ _0923_ _0860_ _0924_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o22ai_1
X_1207_ fifo_dfifo__reg_o7_c_o2_c VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__inv_2
X_1208_ _0927_ _0923_ _0863_ _0924_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__o22ai_1
X_1209_ fifo_dfifo__reg_o7_c_o1_c VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__inv_2
X_1210_ _0928_ _0923_ _0866_ _0924_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o22ai_1
X_1211_ fifo_dfifo__reg_o7_c_o0_c VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__inv_2
X_1212_ _0929_ _0906_ _0869_ _0905_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__o22ai_1
X_1213_ _0785_ _0807_ fifo_dwrite__ptr_o1_c VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__or3_1
X_1214_ _0902_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__or2_4
X_1215_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__clkbuf_2
X_1216_ _0931_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__inv_2
X_1217_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_2
X_1218_ _0896_ _0932_ fifo_dfifo__reg_o6_c_o15_c _0875_ _0934_ VGND VGND VPWR VPWR _0402_
+ sky130_fd_sc_hd__a32o_1
X_1219_ _0895_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__buf_2
X_1220_ _0935_ _0932_ fifo_dfifo__reg_o6_c_o14_c _0878_ _0934_ VGND VGND VPWR VPWR _0401_
+ sky130_fd_sc_hd__a32o_1
X_1221_ _0935_ _0932_ fifo_dfifo__reg_o6_c_o13_c _0880_ _0934_ VGND VGND VPWR VPWR _0400_
+ sky130_fd_sc_hd__a32o_1
X_1222_ _0935_ _0932_ fifo_dfifo__reg_o6_c_o12_c _0881_ _0934_ VGND VGND VPWR VPWR _0399_
+ sky130_fd_sc_hd__a32o_1
X_1223_ _0935_ _0932_ fifo_dfifo__reg_o6_c_o11_c _0882_ _0934_ VGND VGND VPWR VPWR _0398_
+ sky130_fd_sc_hd__a32o_1
X_1224_ _0931_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1225_ _0933_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1226_ _0935_ _0936_ fifo_dfifo__reg_o6_c_o10_c _0884_ _0937_ VGND VGND VPWR VPWR _0397_
+ sky130_fd_sc_hd__a32o_1
X_1227_ _0895_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__buf_2
X_1228_ _0938_ _0936_ fifo_dfifo__reg_o6_c_o9_c _0886_ _0937_ VGND VGND VPWR VPWR _0396_
+ sky130_fd_sc_hd__a32o_1
X_1229_ _0938_ _0936_ fifo_dfifo__reg_o6_c_o8_c _0888_ _0937_ VGND VGND VPWR VPWR _0395_
+ sky130_fd_sc_hd__a32o_1
X_1230_ _0938_ _0936_ fifo_dfifo__reg_o6_c_o7_c _0889_ _0937_ VGND VGND VPWR VPWR _0394_
+ sky130_fd_sc_hd__a32o_1
X_1231_ _0938_ _0936_ fifo_dfifo__reg_o6_c_o6_c _0890_ _0937_ VGND VGND VPWR VPWR _0393_
+ sky130_fd_sc_hd__a32o_1
X_1232_ _0931_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1233_ _0933_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1234_ _0938_ _0939_ fifo_dfifo__reg_o6_c_o5_c _0892_ _0940_ VGND VGND VPWR VPWR _0392_
+ sky130_fd_sc_hd__a32o_1
X_1235_ _0895_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__buf_2
X_1236_ _0941_ _0939_ fifo_dfifo__reg_o6_c_o4_c _0894_ _0940_ VGND VGND VPWR VPWR _0391_
+ sky130_fd_sc_hd__a32o_1
X_1237_ _0941_ _0939_ fifo_dfifo__reg_o6_c_o3_c _0897_ _0940_ VGND VGND VPWR VPWR _0390_
+ sky130_fd_sc_hd__a32o_1
X_1238_ _0941_ _0939_ fifo_dfifo__reg_o6_c_o2_c _0898_ _0940_ VGND VGND VPWR VPWR _0389_
+ sky130_fd_sc_hd__a32o_1
X_1239_ _0941_ _0939_ fifo_dfifo__reg_o6_c_o1_c _0899_ _0940_ VGND VGND VPWR VPWR _0388_
+ sky130_fd_sc_hd__a32o_1
X_1240_ _0941_ _0931_ fifo_dfifo__reg_o6_c_o0_c _0900_ _0933_ VGND VGND VPWR VPWR _0387_
+ sky130_fd_sc_hd__a32o_1
X_1241_ fifo_dfifo__reg_o5_c_o15_c VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__inv_2
X_1242_ _0782_ _0783_ _0902_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__or3_4
X_1243_ _0781_ _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__nand2_4
X_1244_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__clkbuf_2
X_1245_ _0943_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__clkbuf_2
X_1246_ _0942_ _0945_ _0909_ _0946_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o22ai_1
X_1247_ fifo_dfifo__reg_o5_c_o14_c VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__inv_2
X_1248_ _0947_ _0945_ _0819_ _0946_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o22ai_1
X_1249_ fifo_dfifo__reg_o5_c_o13_c VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__inv_2
X_1250_ _0948_ _0945_ _0822_ _0946_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__o22ai_1
X_1251_ fifo_dfifo__reg_o5_c_o12_c VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__inv_2
X_1252_ _0949_ _0945_ _0826_ _0946_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o22ai_1
X_1253_ fifo_dfifo__reg_o5_c_o11_c VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__inv_2
X_1254_ _0950_ _0945_ _0830_ _0946_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o22ai_1
X_1255_ fifo_dfifo__reg_o5_c_o10_c VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__inv_2
X_1256_ _0944_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__clkbuf_2
X_1257_ _0943_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__clkbuf_2
X_1258_ _0951_ _0952_ _0833_ _0953_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o22ai_1
X_1259_ fifo_dfifo__reg_o5_c_o9_c VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__inv_2
X_1260_ _0954_ _0952_ _0838_ _0953_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__o22ai_1
X_1261_ fifo_dfifo__reg_o5_c_o8_c VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__inv_2
X_1262_ _0955_ _0952_ _0841_ _0953_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o22ai_1
X_1263_ fifo_dfifo__reg_o5_c_o7_c VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__inv_2
X_1264_ _0956_ _0952_ _0845_ _0953_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__o22ai_1
X_1265_ fifo_dfifo__reg_o5_c_o6_c VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__inv_2
X_1266_ _0957_ _0952_ _0849_ _0953_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__o22ai_1
X_1267_ fifo_dfifo__reg_o5_c_o5_c VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__inv_2
X_1268_ _0944_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__clkbuf_2
X_1269_ _0943_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__clkbuf_2
X_1270_ _0958_ _0959_ _0852_ _0960_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__o22ai_1
X_1271_ fifo_dfifo__reg_o5_c_o4_c VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__inv_2
X_1272_ _0961_ _0959_ _0857_ _0960_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__o22ai_1
X_1273_ fifo_dfifo__reg_o5_c_o3_c VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__inv_2
X_1274_ _0962_ _0959_ _0860_ _0960_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o22ai_1
X_1275_ fifo_dfifo__reg_o5_c_o2_c VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__inv_2
X_1276_ _0963_ _0959_ _0863_ _0960_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__o22ai_1
X_1277_ fifo_dfifo__reg_o5_c_o1_c VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__inv_2
X_1278_ _0964_ _0959_ _0866_ _0960_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__o22ai_1
X_1279_ fifo_dfifo__reg_o5_c_o0_c VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__inv_2
X_1280_ _0965_ _0944_ _0869_ _0943_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o22ai_1
X_1281_ fifo_dfifo__reg_o4_c_o15_c VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__inv_2
X_1282_ _0792_ _0902_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__or2_4
X_1283_ _0781_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__nand2_4
X_1284_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__buf_2
X_1285_ _0967_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__clkbuf_2
X_1286_ _0966_ _0969_ _0909_ _0970_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__o22ai_1
X_1287_ fifo_dfifo__reg_o4_c_o14_c VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__inv_2
X_1288_ _0971_ _0969_ _0819_ _0970_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o22ai_1
X_1289_ fifo_dfifo__reg_o4_c_o13_c VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__inv_2
X_1290_ _0972_ _0969_ _0822_ _0970_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o22ai_1
X_1291_ fifo_dfifo__reg_o4_c_o12_c VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__inv_2
X_1292_ _0973_ _0969_ _0826_ _0970_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o22ai_1
X_1293_ fifo_dfifo__reg_o4_c_o11_c VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__inv_2
X_1294_ _0974_ _0969_ _0830_ _0970_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o22ai_1
X_1295_ fifo_dfifo__reg_o4_c_o10_c VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__inv_2
X_1296_ _0968_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__clkbuf_2
X_1297_ _0967_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__clkbuf_2
X_1298_ _0975_ _0976_ _0833_ _0977_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o22ai_1
X_1299_ fifo_dfifo__reg_o4_c_o9_c VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__inv_2
X_1300_ _0978_ _0976_ _0838_ _0977_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o22ai_1
X_1301_ fifo_dfifo__reg_o4_c_o8_c VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__inv_2
X_1302_ _0979_ _0976_ _0841_ _0977_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__o22ai_1
X_1303_ fifo_dfifo__reg_o4_c_o7_c VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__inv_2
X_1304_ _0980_ _0976_ _0845_ _0977_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o22ai_1
X_1305_ fifo_dfifo__reg_o4_c_o6_c VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__inv_2
X_1306_ _0981_ _0976_ _0849_ _0977_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o22ai_1
X_1307_ fifo_dfifo__reg_o4_c_o5_c VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__inv_2
X_1308_ _0968_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__clkbuf_2
X_1309_ _0967_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__clkbuf_2
X_1310_ _0982_ _0983_ _0852_ _0984_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__o22ai_1
X_1311_ fifo_dfifo__reg_o4_c_o4_c VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__inv_2
X_1312_ _0985_ _0983_ _0857_ _0984_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__o22ai_1
X_1313_ fifo_dfifo__reg_o4_c_o3_c VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__inv_2
X_1314_ _0986_ _0983_ _0860_ _0984_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o22ai_1
X_1315_ fifo_dfifo__reg_o4_c_o2_c VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__inv_2
X_1316_ _0987_ _0983_ _0863_ _0984_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o22ai_1
X_1317_ fifo_dfifo__reg_o4_c_o1_c VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__inv_2
X_1318_ _0988_ _0983_ _0866_ _0984_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__o22ai_1
X_1319_ fifo_dfifo__reg_o4_c_o0_c VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__inv_2
X_1320_ _0989_ _0968_ _0869_ _0967_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o22ai_1
X_1321_ fifo_dfifo__reg_o3_c_o15_c VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__inv_2
X_1322_ _0796_ _0808_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__or2_1
X_1323_ _0904_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__or2_4
X_1324_ _0781_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__nand2_4
X_1325_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__clkbuf_2
X_1326_ _0992_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__clkbuf_2
X_1327_ _0990_ _0994_ _0909_ _0995_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o22ai_1
X_1328_ fifo_dfifo__reg_o3_c_o14_c VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__inv_2
X_1329_ _0996_ _0994_ _0819_ _0995_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o22ai_1
X_1330_ fifo_dfifo__reg_o3_c_o13_c VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__inv_2
X_1331_ _0997_ _0994_ _0822_ _0995_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o22ai_1
X_1332_ fifo_dfifo__reg_o3_c_o12_c VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__inv_2
X_1333_ _0998_ _0994_ _0826_ _0995_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o22ai_1
X_1334_ fifo_dfifo__reg_o3_c_o11_c VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__inv_2
X_1335_ _0999_ _0994_ _0830_ _0995_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o22ai_1
X_1336_ fifo_dfifo__reg_o3_c_o10_c VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
X_1337_ _0993_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_2
X_1338_ _0992_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__clkbuf_2
X_1339_ _1000_ _1001_ _0833_ _1002_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__o22ai_1
X_1340_ fifo_dfifo__reg_o3_c_o9_c VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__inv_2
X_1341_ _1003_ _1001_ _0838_ _1002_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o22ai_1
X_1342_ fifo_dfifo__reg_o3_c_o8_c VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__inv_2
X_1343_ _1004_ _1001_ _0841_ _1002_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o22ai_1
X_1344_ fifo_dfifo__reg_o3_c_o7_c VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__inv_2
X_1345_ _1005_ _1001_ _0845_ _1002_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o22ai_1
X_1346_ fifo_dfifo__reg_o3_c_o6_c VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__inv_2
X_1347_ _1006_ _1001_ _0849_ _1002_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o22ai_1
X_1348_ fifo_dfifo__reg_o3_c_o5_c VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__inv_2
X_1349_ _0993_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1350_ _0992_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1351_ _1007_ _1008_ _0852_ _1009_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o22ai_1
X_1352_ fifo_dfifo__reg_o3_c_o4_c VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__inv_2
X_1353_ _1010_ _1008_ _0857_ _1009_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o22ai_1
X_1354_ fifo_dfifo__reg_o3_c_o3_c VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__inv_2
X_1355_ _0451_ _1008_ _0860_ _1009_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o22ai_1
X_1356_ fifo_dfifo__reg_o3_c_o2_c VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__inv_2
X_1357_ _0452_ _1008_ _0863_ _1009_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o22ai_1
X_1358_ fifo_dfifo__reg_o3_c_o1_c VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__inv_2
X_1359_ _0453_ _1008_ _0866_ _1009_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o22ai_1
X_1360_ fifo_dfifo__reg_o3_c_o0_c VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__inv_2
X_1361_ _0454_ _0993_ _0869_ _0992_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__o22ai_1
X_1362_ _0895_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_2
X_1363_ _0930_ _0991_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or2_4
X_1364_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_2
X_1365_ _0456_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__inv_2
X_1366_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_2
X_1367_ _0455_ _0457_ fifo_dfifo__reg_o2_c_o15_c _0875_ _0459_ VGND VGND VPWR VPWR _0338_
+ sky130_fd_sc_hd__a32o_1
X_1368_ _0455_ _0457_ fifo_dfifo__reg_o2_c_o14_c _0878_ _0459_ VGND VGND VPWR VPWR _0337_
+ sky130_fd_sc_hd__a32o_1
X_1369_ _0455_ _0457_ fifo_dfifo__reg_o2_c_o13_c _0880_ _0459_ VGND VGND VPWR VPWR _0336_
+ sky130_fd_sc_hd__a32o_1
X_1370_ _0455_ _0457_ fifo_dfifo__reg_o2_c_o12_c _0881_ _0459_ VGND VGND VPWR VPWR _0335_
+ sky130_fd_sc_hd__a32o_1
X_1371_ _0455_ _0457_ fifo_dfifo__reg_o2_c_o11_c _0882_ _0459_ VGND VGND VPWR VPWR _0334_
+ sky130_fd_sc_hd__a32o_1
X_1372_ _0780_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_4
X_1373_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1374_ _0456_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1375_ _0458_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1376_ _0461_ _0462_ fifo_dfifo__reg_o2_c_o10_c _0884_ _0463_ VGND VGND VPWR VPWR _0333_
+ sky130_fd_sc_hd__a32o_1
X_1377_ _0461_ _0462_ fifo_dfifo__reg_o2_c_o9_c _0886_ _0463_ VGND VGND VPWR VPWR _0332_
+ sky130_fd_sc_hd__a32o_1
X_1378_ _0461_ _0462_ fifo_dfifo__reg_o2_c_o8_c _0888_ _0463_ VGND VGND VPWR VPWR _0331_
+ sky130_fd_sc_hd__a32o_1
X_1379_ _0461_ _0462_ fifo_dfifo__reg_o2_c_o7_c _0889_ _0463_ VGND VGND VPWR VPWR _0330_
+ sky130_fd_sc_hd__a32o_1
X_1380_ _0461_ _0462_ fifo_dfifo__reg_o2_c_o6_c _0890_ _0463_ VGND VGND VPWR VPWR _0329_
+ sky130_fd_sc_hd__a32o_1
X_1381_ _0460_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1382_ _0456_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1383_ _0458_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1384_ _0464_ _0465_ fifo_dfifo__reg_o2_c_o5_c _0892_ _0466_ VGND VGND VPWR VPWR _0328_
+ sky130_fd_sc_hd__a32o_1
X_1385_ _0464_ _0465_ fifo_dfifo__reg_o2_c_o4_c _0894_ _0466_ VGND VGND VPWR VPWR _0327_
+ sky130_fd_sc_hd__a32o_1
X_1386_ _0464_ _0465_ fifo_dfifo__reg_o2_c_o3_c _0897_ _0466_ VGND VGND VPWR VPWR _0326_
+ sky130_fd_sc_hd__a32o_1
X_1387_ _0464_ _0465_ fifo_dfifo__reg_o2_c_o2_c _0898_ _0466_ VGND VGND VPWR VPWR _0325_
+ sky130_fd_sc_hd__a32o_1
X_1388_ _0464_ _0465_ fifo_dfifo__reg_o2_c_o1_c _0899_ _0466_ VGND VGND VPWR VPWR _0324_
+ sky130_fd_sc_hd__a32o_1
X_1389_ _0460_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_2
X_1390_ _0467_ _0456_ fifo_dfifo__reg_o2_c_o0_c _0900_ _0458_ VGND VGND VPWR VPWR _0323_
+ sky130_fd_sc_hd__a32o_1
X_1391_ fifo_dfifo__reg_o1_c_o15_c VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__inv_2
X_1392_ _0782_ _0783_ _0991_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or3_4
X_1393_ _0870_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nand2_4
X_1394_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_2
X_1395_ _0469_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_2
X_1396_ _0468_ _0471_ _0908_ _0472_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__o22ai_1
X_1397_ fifo_dfifo__reg_o1_c_o14_c VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__inv_2
X_1398_ _0473_ _0471_ _0818_ _0472_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o22ai_1
X_1399_ fifo_dfifo__reg_o1_c_o13_c VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__inv_2
X_1400_ _0474_ _0471_ _0821_ _0472_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__o22ai_1
X_1401_ fifo_dfifo__reg_o1_c_o12_c VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__inv_2
X_1402_ _0475_ _0471_ _0825_ _0472_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o22ai_1
X_1403_ fifo_dfifo__reg_o1_c_o11_c VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__inv_2
X_1404_ _0476_ _0471_ _0829_ _0472_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o22ai_1
X_1405_ fifo_dfifo__reg_o1_c_o10_c VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__inv_2
X_1406_ _0470_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_2
X_1407_ _0469_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_2
X_1408_ _0477_ _0478_ _0832_ _0479_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o22ai_1
X_1409_ fifo_dfifo__reg_o1_c_o9_c VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__inv_2
X_1410_ _0480_ _0478_ _0837_ _0479_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o22ai_1
X_1411_ fifo_dfifo__reg_o1_c_o8_c VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__inv_2
X_1412_ _0481_ _0478_ _0840_ _0479_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o22ai_1
X_1413_ fifo_dfifo__reg_o1_c_o7_c VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__inv_2
X_1414_ _0482_ _0478_ _0844_ _0479_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__o22ai_1
X_1415_ fifo_dfifo__reg_o1_c_o6_c VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__inv_2
X_1416_ _0483_ _0478_ _0848_ _0479_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__o22ai_1
X_1417_ fifo_dfifo__reg_o1_c_o5_c VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__inv_2
X_1418_ _0470_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__clkbuf_2
X_1419_ _0469_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__clkbuf_2
X_1420_ _0484_ _0485_ _0851_ _0486_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__o22ai_1
X_1421_ fifo_dfifo__reg_o1_c_o4_c VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__inv_2
X_1422_ _0487_ _0485_ _0856_ _0486_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__o22ai_1
X_1423_ fifo_dfifo__reg_o1_c_o3_c VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__inv_2
X_1424_ _0488_ _0485_ _0859_ _0486_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__o22ai_1
X_1425_ fifo_dfifo__reg_o1_c_o2_c VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__inv_2
X_1426_ _0489_ _0485_ _0862_ _0486_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o22ai_1
X_1427_ fifo_dfifo__reg_o1_c_o1_c VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__inv_2
X_1428_ _0490_ _0485_ _0865_ _0486_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o22ai_1
X_1429_ fifo_dfifo__reg_o1_c_o0_c VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__inv_2
X_1430_ _0491_ _0470_ _0868_ _0469_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__o22ai_1
X_1431_ _0796_ _0903_ _0808_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o21ai_2
X_1432_ _0930_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or2_2
X_1433_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__clkbuf_2
X_1434_ _0493_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__inv_2
X_1435_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_2
X_1436_ _0467_ _0494_ fifo_dfifo__reg_o14_c_o15_c _0875_ _0496_ VGND VGND VPWR VPWR _0306_
+ sky130_fd_sc_hd__a32o_1
X_1437_ _0467_ _0494_ fifo_dfifo__reg_o14_c_o14_c _0878_ _0496_ VGND VGND VPWR VPWR _0305_
+ sky130_fd_sc_hd__a32o_1
X_1438_ _0467_ _0494_ fifo_dfifo__reg_o14_c_o13_c _0880_ _0496_ VGND VGND VPWR VPWR _0304_
+ sky130_fd_sc_hd__a32o_1
X_1439_ _0467_ _0494_ fifo_dfifo__reg_o14_c_o12_c _0881_ _0496_ VGND VGND VPWR VPWR _0303_
+ sky130_fd_sc_hd__a32o_1
X_1440_ _0460_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_2
X_1441_ _0497_ _0494_ fifo_dfifo__reg_o14_c_o11_c _0882_ _0496_ VGND VGND VPWR VPWR _0302_
+ sky130_fd_sc_hd__a32o_1
X_1442_ _0493_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__clkbuf_2
X_1443_ _0495_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_2
X_1444_ _0497_ _0498_ fifo_dfifo__reg_o14_c_o10_c _0884_ _0499_ VGND VGND VPWR VPWR _0301_
+ sky130_fd_sc_hd__a32o_1
X_1445_ _0497_ _0498_ fifo_dfifo__reg_o14_c_o9_c _0886_ _0499_ VGND VGND VPWR VPWR _0300_
+ sky130_fd_sc_hd__a32o_1
X_1446_ _0497_ _0498_ fifo_dfifo__reg_o14_c_o8_c _0888_ _0499_ VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__a32o_1
X_1447_ _0497_ _0498_ fifo_dfifo__reg_o14_c_o7_c _0889_ _0499_ VGND VGND VPWR VPWR _0298_
+ sky130_fd_sc_hd__a32o_1
X_1448_ _0460_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_2
X_1449_ _0500_ _0498_ fifo_dfifo__reg_o14_c_o6_c _0890_ _0499_ VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__a32o_1
X_1450_ _0493_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1451_ _0495_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1452_ _0500_ _0501_ fifo_dfifo__reg_o14_c_o5_c _0892_ _0502_ VGND VGND VPWR VPWR _0296_
+ sky130_fd_sc_hd__a32o_1
X_1453_ _0500_ _0501_ fifo_dfifo__reg_o14_c_o4_c _0894_ _0502_ VGND VGND VPWR VPWR _0295_
+ sky130_fd_sc_hd__a32o_1
X_1454_ _0500_ _0501_ fifo_dfifo__reg_o14_c_o3_c _0897_ _0502_ VGND VGND VPWR VPWR _0294_
+ sky130_fd_sc_hd__a32o_1
X_1455_ _0500_ _0501_ fifo_dfifo__reg_o14_c_o2_c _0898_ _0502_ VGND VGND VPWR VPWR _0293_
+ sky130_fd_sc_hd__a32o_1
X_1456_ _0780_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1457_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_2
X_1458_ _0504_ _0501_ fifo_dfifo__reg_o14_c_o1_c _0899_ _0502_ VGND VGND VPWR VPWR _0292_
+ sky130_fd_sc_hd__a32o_1
X_1459_ _0504_ _0493_ fifo_dfifo__reg_o14_c_o0_c _0900_ _0495_ VGND VGND VPWR VPWR _0291_
+ sky130_fd_sc_hd__a32o_1
X_1460_ _0782_ _0783_ _0903_ _0492_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__or4_4
X_1461_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1462_ _0505_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__clkinv_2
X_1463_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__clkbuf_2
X_1464_ _0504_ _0506_ fifo_dfifo__reg_o13_c_o15_c _0875_ _0508_ VGND VGND VPWR VPWR _0290_
+ sky130_fd_sc_hd__a32o_1
X_1465_ _0504_ _0506_ fifo_dfifo__reg_o13_c_o14_c _0878_ _0508_ VGND VGND VPWR VPWR _0289_
+ sky130_fd_sc_hd__a32o_1
X_1466_ _0504_ _0506_ fifo_dfifo__reg_o13_c_o13_c _0880_ _0508_ VGND VGND VPWR VPWR _0288_
+ sky130_fd_sc_hd__a32o_1
X_1467_ _0503_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_2
X_1468_ _0509_ _0506_ fifo_dfifo__reg_o13_c_o12_c _0881_ _0508_ VGND VGND VPWR VPWR _0287_
+ sky130_fd_sc_hd__a32o_1
X_1469_ _0509_ _0506_ fifo_dfifo__reg_o13_c_o11_c _0882_ _0508_ VGND VGND VPWR VPWR _0286_
+ sky130_fd_sc_hd__a32o_1
X_1470_ _0505_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_2
X_1471_ _0507_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_2
X_1472_ _0509_ _0510_ fifo_dfifo__reg_o13_c_o10_c _0884_ _0511_ VGND VGND VPWR VPWR _0285_
+ sky130_fd_sc_hd__a32o_1
X_1473_ _0509_ _0510_ fifo_dfifo__reg_o13_c_o9_c _0886_ _0511_ VGND VGND VPWR VPWR _0284_
+ sky130_fd_sc_hd__a32o_1
X_1474_ _0509_ _0510_ fifo_dfifo__reg_o13_c_o8_c _0888_ _0511_ VGND VGND VPWR VPWR _0283_
+ sky130_fd_sc_hd__a32o_1
X_1475_ _0503_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__buf_2
X_1476_ _0512_ _0510_ fifo_dfifo__reg_o13_c_o7_c _0889_ _0511_ VGND VGND VPWR VPWR _0282_
+ sky130_fd_sc_hd__a32o_1
X_1477_ _0512_ _0510_ fifo_dfifo__reg_o13_c_o6_c _0890_ _0511_ VGND VGND VPWR VPWR _0281_
+ sky130_fd_sc_hd__a32o_1
X_1478_ _0505_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1479_ _0507_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1480_ _0512_ _0513_ fifo_dfifo__reg_o13_c_o5_c _0892_ _0514_ VGND VGND VPWR VPWR _0280_
+ sky130_fd_sc_hd__a32o_1
X_1481_ _0512_ _0513_ fifo_dfifo__reg_o13_c_o4_c _0894_ _0514_ VGND VGND VPWR VPWR _0279_
+ sky130_fd_sc_hd__a32o_1
X_1482_ _0512_ _0513_ fifo_dfifo__reg_o13_c_o3_c _0897_ _0514_ VGND VGND VPWR VPWR _0278_
+ sky130_fd_sc_hd__a32o_1
X_1483_ _0503_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__buf_2
X_1484_ _0515_ _0513_ fifo_dfifo__reg_o13_c_o2_c _0898_ _0514_ VGND VGND VPWR VPWR _0277_
+ sky130_fd_sc_hd__a32o_1
X_1485_ _0515_ _0513_ fifo_dfifo__reg_o13_c_o1_c _0899_ _0514_ VGND VGND VPWR VPWR _0276_
+ sky130_fd_sc_hd__a32o_1
X_1486_ _0515_ _0505_ fifo_dfifo__reg_o13_c_o0_c _0900_ _0507_ VGND VGND VPWR VPWR _0275_
+ sky130_fd_sc_hd__a32o_1
X_1487_ _0792_ _0903_ _0492_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__or3_4
X_1488_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1489_ _0516_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__clkinv_2
X_1490_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1491_ _0515_ _0517_ fifo_dfifo__reg_o12_c_o15_c net7 _0519_ VGND VGND VPWR VPWR _0274_
+ sky130_fd_sc_hd__a32o_1
X_1492_ _0515_ _0517_ fifo_dfifo__reg_o12_c_o14_c net6 _0519_ VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__a32o_1
X_1493_ _0503_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_2
X_1494_ _0520_ _0517_ fifo_dfifo__reg_o12_c_o13_c net5 _0519_ VGND VGND VPWR VPWR _0272_
+ sky130_fd_sc_hd__a32o_1
X_1495_ _0520_ _0517_ fifo_dfifo__reg_o12_c_o12_c net4 _0519_ VGND VGND VPWR VPWR _0271_
+ sky130_fd_sc_hd__a32o_1
X_1496_ _0520_ _0517_ fifo_dfifo__reg_o12_c_o11_c net3 _0519_ VGND VGND VPWR VPWR _0270_
+ sky130_fd_sc_hd__a32o_1
X_1497_ _0516_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_2
X_1498_ _0518_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_2
X_1499_ _0520_ _0521_ fifo_dfifo__reg_o12_c_o10_c net2 _0522_ VGND VGND VPWR VPWR _0269_
+ sky130_fd_sc_hd__a32o_1
X_1500_ _0520_ _0521_ fifo_dfifo__reg_o12_c_o9_c net16 _0522_ VGND VGND VPWR VPWR _0268_
+ sky130_fd_sc_hd__a32o_1
X_1501_ _0780_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1502_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_2
X_1503_ _0524_ _0521_ fifo_dfifo__reg_o12_c_o8_c net15 _0522_ VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__a32o_1
X_1504_ _0524_ _0521_ fifo_dfifo__reg_o12_c_o7_c net14 _0522_ VGND VGND VPWR VPWR _0266_
+ sky130_fd_sc_hd__a32o_1
X_1505_ _0524_ _0521_ fifo_dfifo__reg_o12_c_o6_c net13 _0522_ VGND VGND VPWR VPWR _0265_
+ sky130_fd_sc_hd__a32o_1
X_1506_ _0516_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_2
X_1507_ _0518_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1508_ _0524_ _0525_ fifo_dfifo__reg_o12_c_o5_c net12 _0526_ VGND VGND VPWR VPWR _0264_
+ sky130_fd_sc_hd__a32o_1
X_1509_ _0524_ _0525_ fifo_dfifo__reg_o12_c_o4_c net11 _0526_ VGND VGND VPWR VPWR _0263_
+ sky130_fd_sc_hd__a32o_1
X_1510_ _0523_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__buf_2
X_1511_ _0527_ _0525_ fifo_dfifo__reg_o12_c_o3_c net10 _0526_ VGND VGND VPWR VPWR _0262_
+ sky130_fd_sc_hd__a32o_1
X_1512_ _0527_ _0525_ fifo_dfifo__reg_o12_c_o2_c net9 _0526_ VGND VGND VPWR VPWR _0261_
+ sky130_fd_sc_hd__a32o_1
X_1513_ _0527_ _0525_ fifo_dfifo__reg_o12_c_o1_c net8 _0526_ VGND VGND VPWR VPWR _0260_
+ sky130_fd_sc_hd__a32o_1
X_1514_ _0527_ _0516_ fifo_dfifo__reg_o12_c_o0_c net1 _0518_ VGND VGND VPWR VPWR _0259_
+ sky130_fd_sc_hd__a32o_1
X_1515_ fifo_dfifo__reg_o11_c_o15_c VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__inv_2
X_1516_ _0809_ _0904_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or2_4
X_1517_ _0870_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nand2_2
X_1518_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__clkbuf_2
X_1519_ _0529_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__clkbuf_2
X_1520_ _0528_ _0531_ _0908_ _0532_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__o22ai_1
X_1521_ fifo_dfifo__reg_o11_c_o14_c VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__inv_2
X_1522_ _0533_ _0531_ _0818_ _0532_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__o22ai_1
X_1523_ fifo_dfifo__reg_o11_c_o13_c VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__inv_2
X_1524_ _0534_ _0531_ _0821_ _0532_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o22ai_1
X_1525_ fifo_dfifo__reg_o11_c_o12_c VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__inv_2
X_1526_ _0535_ _0531_ _0825_ _0532_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__o22ai_1
X_1527_ fifo_dfifo__reg_o11_c_o11_c VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__inv_2
X_1528_ _0536_ _0531_ _0829_ _0532_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__o22ai_1
X_1529_ fifo_dfifo__reg_o11_c_o10_c VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__inv_2
X_1530_ _0530_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__buf_2
X_1531_ _0529_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__buf_2
X_1532_ _0537_ _0538_ _0832_ _0539_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__o22ai_1
X_1533_ fifo_dfifo__reg_o11_c_o9_c VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__inv_2
X_1534_ _0540_ _0538_ _0837_ _0539_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__o22ai_1
X_1535_ fifo_dfifo__reg_o11_c_o8_c VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__inv_2
X_1536_ _0541_ _0538_ _0840_ _0539_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o22ai_1
X_1537_ fifo_dfifo__reg_o11_c_o7_c VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__inv_2
X_1538_ _0542_ _0538_ _0844_ _0539_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__o22ai_1
X_1539_ fifo_dfifo__reg_o11_c_o6_c VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__inv_2
X_1540_ _0543_ _0538_ _0848_ _0539_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o22ai_1
X_1541_ fifo_dfifo__reg_o11_c_o5_c VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__inv_2
X_1542_ _0530_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__clkbuf_2
X_1543_ _0529_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_2
X_1544_ _0544_ _0545_ _0851_ _0546_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o22ai_1
X_1545_ fifo_dfifo__reg_o11_c_o4_c VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__inv_2
X_1546_ _0547_ _0545_ _0856_ _0546_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o22ai_1
X_1547_ fifo_dfifo__reg_o11_c_o3_c VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__inv_2
X_1548_ _0548_ _0545_ _0859_ _0546_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o22ai_1
X_1549_ fifo_dfifo__reg_o11_c_o2_c VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__inv_2
X_1550_ _0549_ _0545_ _0862_ _0546_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o22ai_1
X_1551_ fifo_dfifo__reg_o11_c_o1_c VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__inv_2
X_1552_ _0550_ _0545_ _0865_ _0546_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o22ai_1
X_1553_ fifo_dfifo__reg_o11_c_o0_c VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__inv_2
X_1554_ _0551_ _0530_ _0868_ _0529_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__o22ai_1
X_1555_ _0809_ _0930_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or2_2
X_1556_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_2
X_1557_ _0552_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__inv_2
X_1558_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_2
X_1559_ _0527_ _0553_ fifo_dfifo__reg_o10_c_o15_c net7 _0555_ VGND VGND VPWR VPWR _0242_
+ sky130_fd_sc_hd__a32o_1
X_1560_ _0523_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__clkbuf_2
X_1561_ _0556_ _0553_ fifo_dfifo__reg_o10_c_o14_c net6 _0555_ VGND VGND VPWR VPWR _0241_
+ sky130_fd_sc_hd__a32o_1
X_1562_ _0556_ _0553_ fifo_dfifo__reg_o10_c_o13_c net5 _0555_ VGND VGND VPWR VPWR _0240_
+ sky130_fd_sc_hd__a32o_1
X_1563_ _0556_ _0553_ fifo_dfifo__reg_o10_c_o12_c net4 _0555_ VGND VGND VPWR VPWR _0239_
+ sky130_fd_sc_hd__a32o_1
X_1564_ _0556_ _0553_ fifo_dfifo__reg_o10_c_o11_c net3 _0555_ VGND VGND VPWR VPWR _0238_
+ sky130_fd_sc_hd__a32o_1
X_1565_ _0552_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__clkbuf_2
X_1566_ _0554_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_2
X_1567_ _0556_ _0557_ fifo_dfifo__reg_o10_c_o10_c net2 _0558_ VGND VGND VPWR VPWR _0237_
+ sky130_fd_sc_hd__a32o_1
X_1568_ _0523_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__buf_2
X_1569_ _0559_ _0557_ fifo_dfifo__reg_o10_c_o9_c net16 _0558_ VGND VGND VPWR VPWR _0236_
+ sky130_fd_sc_hd__a32o_1
X_1570_ _0559_ _0557_ fifo_dfifo__reg_o10_c_o8_c net15 _0558_ VGND VGND VPWR VPWR _0235_
+ sky130_fd_sc_hd__a32o_1
X_1571_ _0559_ _0557_ fifo_dfifo__reg_o10_c_o7_c net14 _0558_ VGND VGND VPWR VPWR _0234_
+ sky130_fd_sc_hd__a32o_1
X_1572_ _0559_ _0557_ fifo_dfifo__reg_o10_c_o6_c net13 _0558_ VGND VGND VPWR VPWR _0233_
+ sky130_fd_sc_hd__a32o_1
X_1573_ _0552_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__clkbuf_2
X_1574_ _0554_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_2
X_1575_ _0559_ _0560_ fifo_dfifo__reg_o10_c_o5_c net12 _0561_ VGND VGND VPWR VPWR _0232_
+ sky130_fd_sc_hd__a32o_1
X_1576_ _0523_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_2
X_1577_ _0562_ _0560_ fifo_dfifo__reg_o10_c_o4_c net11 _0561_ VGND VGND VPWR VPWR _0231_
+ sky130_fd_sc_hd__a32o_1
X_1578_ _0562_ _0560_ fifo_dfifo__reg_o10_c_o3_c net10 _0561_ VGND VGND VPWR VPWR _0230_
+ sky130_fd_sc_hd__a32o_1
X_1579_ _0562_ _0560_ fifo_dfifo__reg_o10_c_o2_c net9 _0561_ VGND VGND VPWR VPWR _0229_
+ sky130_fd_sc_hd__a32o_1
X_1580_ _0562_ _0560_ fifo_dfifo__reg_o10_c_o1_c net8 _0561_ VGND VGND VPWR VPWR _0228_
+ sky130_fd_sc_hd__a32o_1
X_1581_ _0562_ _0552_ fifo_dfifo__reg_o10_c_o0_c net1 _0554_ VGND VGND VPWR VPWR _0227_
+ sky130_fd_sc_hd__a32o_1
X_1582_ _0780_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__buf_4
X_1583_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1584_ _0792_ _0991_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__or2_4
X_1585_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__clkbuf_2
X_1586_ _0565_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__inv_2
X_1587_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_2
X_1588_ _0564_ _0566_ fifo_dfifo__reg_o0_c_o15_c net7 _0568_ VGND VGND VPWR VPWR _0226_
+ sky130_fd_sc_hd__a32o_1
X_1589_ _0564_ _0566_ fifo_dfifo__reg_o0_c_o14_c net6 _0568_ VGND VGND VPWR VPWR _0225_
+ sky130_fd_sc_hd__a32o_1
X_1590_ _0564_ _0566_ fifo_dfifo__reg_o0_c_o13_c net5 _0568_ VGND VGND VPWR VPWR _0224_
+ sky130_fd_sc_hd__a32o_1
X_1591_ _0564_ _0566_ fifo_dfifo__reg_o0_c_o12_c net4 _0568_ VGND VGND VPWR VPWR _0223_
+ sky130_fd_sc_hd__a32o_1
X_1592_ _0564_ _0566_ fifo_dfifo__reg_o0_c_o11_c net3 _0568_ VGND VGND VPWR VPWR _0222_
+ sky130_fd_sc_hd__a32o_1
X_1593_ _0563_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__clkbuf_2
X_1594_ _0565_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_2
X_1595_ _0567_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__clkbuf_2
X_1596_ _0569_ _0570_ fifo_dfifo__reg_o0_c_o10_c net2 _0571_ VGND VGND VPWR VPWR _0221_
+ sky130_fd_sc_hd__a32o_1
X_1597_ _0569_ _0570_ fifo_dfifo__reg_o0_c_o9_c net16 _0571_ VGND VGND VPWR VPWR _0220_
+ sky130_fd_sc_hd__a32o_1
X_1598_ _0569_ _0570_ fifo_dfifo__reg_o0_c_o8_c net15 _0571_ VGND VGND VPWR VPWR _0219_
+ sky130_fd_sc_hd__a32o_1
X_1599_ _0569_ _0570_ fifo_dfifo__reg_o0_c_o7_c net14 _0571_ VGND VGND VPWR VPWR _0218_
+ sky130_fd_sc_hd__a32o_1
X_1600_ _0569_ _0570_ fifo_dfifo__reg_o0_c_o6_c net13 _0571_ VGND VGND VPWR VPWR _0217_
+ sky130_fd_sc_hd__a32o_1
X_1601_ _0563_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1602_ _0565_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1603_ _0567_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1604_ _0572_ _0573_ fifo_dfifo__reg_o0_c_o5_c net12 _0574_ VGND VGND VPWR VPWR _0216_
+ sky130_fd_sc_hd__a32o_1
X_1605_ _0572_ _0573_ fifo_dfifo__reg_o0_c_o4_c net11 _0574_ VGND VGND VPWR VPWR _0215_
+ sky130_fd_sc_hd__a32o_1
X_1606_ _0572_ _0573_ fifo_dfifo__reg_o0_c_o3_c net10 _0574_ VGND VGND VPWR VPWR _0214_
+ sky130_fd_sc_hd__a32o_1
X_1607_ _0572_ _0573_ fifo_dfifo__reg_o0_c_o2_c net9 _0574_ VGND VGND VPWR VPWR _0213_
+ sky130_fd_sc_hd__a32o_1
X_1608_ _0572_ _0573_ fifo_dfifo__reg_o0_c_o1_c net8 _0574_ VGND VGND VPWR VPWR _0212_
+ sky130_fd_sc_hd__a32o_1
X_1609_ _0563_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_2
X_1610_ _0575_ _0565_ fifo_dfifo__reg_o0_c_o0_c net1 _0567_ VGND VGND VPWR VPWR _0211_
+ sky130_fd_sc_hd__a32o_1
X_1611_ net18 VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__inv_2
X_1612_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__clkbuf_2
X_1613_ dsmod_daccu1_o15_c VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__inv_2
X_1614_ net25 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__inv_2
X_1615_ net22 _0028_ net23 VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__and3_1
X_1616_ _0580_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_1617_ net24 _0141_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nand2_1
X_1618_ _0579_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or2_1
X_1619_ _0578_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nor2_1
X_1620_ _0578_ _0582_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__a21oi_1
X_1621_ net25 VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1622_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1623_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1624_ net23 _0034_ net24 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and3_1
X_1625_ _0588_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1626_ dsmod_daccu1_o14_c VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__inv_2
X_1627_ _0587_ _0154_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nand2_1
X_1628_ _0587_ _0154_ dsmod_daccu1_o14_c _0589_ _0590_ VGND VGND VPWR VPWR _0591_
+ sky130_fd_sc_hd__a32o_1
X_1629_ net24 _0121_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2_1
X_1630_ _0592_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_2
X_1631_ dsmod_daccu1_o13_c VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__inv_2
X_1632_ _0586_ _0151_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nand2_1
X_1633_ _0593_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__and2_1
X_1634_ _0587_ _0151_ dsmod_daccu1_o13_c _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a31o_1
X_1635_ net24 _0046_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__and2_1
X_1636_ _0597_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1637_ dsmod_daccu1_o12_c VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__inv_2
X_1638_ _0586_ _0148_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__nand2_1
X_1639_ _0586_ _0148_ dsmod_daccu1_o12_c _0598_ _0599_ VGND VGND VPWR VPWR _0600_
+ sky130_fd_sc_hd__a32o_1
X_1640_ net25 _0143_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and2_1
X_1641_ dsmod_daccu1_o11_c _0601_ dsmod_daccu1_o11_c _0601_ VGND VGND VPWR VPWR _0602_
+ sky130_fd_sc_hd__o2bb2a_1
X_1642_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__inv_2
X_1643_ _0585_ _0136_ dsmod_daccu1_o10_c VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a21oi_1
X_1644_ _0585_ _0136_ dsmod_daccu1_o10_c _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a31o_1
X_1645_ _0603_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
X_1646_ net25 _0125_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__and2_1
X_1647_ _0585_ _0070_ dsmod_daccu1_o8_c dsmod_daccu1_o9_c _0607_ VGND VGND VPWR VPWR _0608_
+ sky130_fd_sc_hd__a32o_1
X_1648_ dsmod_daccu1_o9_c _0607_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__o21ai_1
X_1649_ dsmod_daccu1_o7_c VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__inv_2
X_1650_ net24 net23 net22 net25 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or4_2
X_1651_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__clkbuf_2
X_1652_ _0159_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nand2_1
X_1653_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__inv_2
X_1654_ _0612_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1655_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1656_ dsmod_daccu1_o7_c _0614_ _0156_ _0616_ dsmod_daccu1_o6_c VGND VGND VPWR VPWR _0617_
+ sky130_fd_sc_hd__o2111ai_1
X_1657_ _0610_ _0613_ dsmod_daccu1_o7_c _0614_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__o22a_1
X_1658_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__inv_2
X_1659_ _0156_ _0615_ dsmod_daccu1_o6_c VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a21oi_1
X_1660_ _0156_ _0616_ dsmod_daccu1_o6_c _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a31o_1
X_1661_ _0619_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or2_1
X_1662_ _0153_ _0615_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__and2_1
X_1663_ _0150_ _0616_ dsmod_daccu1_o4_c dsmod_daccu1_o5_c _0623_ VGND VGND VPWR VPWR _0624_
+ sky130_fd_sc_hd__a32o_1
X_1664_ dsmod_daccu1_o5_c _0623_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__o21ai_1
X_1665_ _0622_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or2_1
X_1666_ dsmod_daccu1_o5_c _0623_ dsmod_daccu1_o5_c _0623_ VGND VGND VPWR VPWR _0627_
+ sky130_fd_sc_hd__o2bb2a_1
X_1667_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__inv_2
X_1668_ _0150_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__inv_2
X_1669_ _0611_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__inv_2
X_1670_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1671_ dsmod_daccu1_o4_c VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__inv_2
X_1672_ _0629_ _0631_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o21a_1
X_1673_ _0150_ _0616_ dsmod_daccu1_o4_c _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a31o_1
X_1674_ _0147_ _0611_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__and2_1
X_1675_ dsmod_daccu1_o3_c _0635_ dsmod_daccu1_o3_c _0635_ VGND VGND VPWR VPWR _0636_
+ sky130_fd_sc_hd__o2bb2a_1
X_1676_ _0140_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__inv_2
X_1677_ dsmod_daccu1_o2_c VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__inv_2
X_1678_ _0637_ _0630_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__o21a_1
X_1679_ _0140_ _0612_ dsmod_daccu1_o2_c _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a31o_1
X_1680_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__inv_2
X_1681_ _0133_ _0611_ dsmod_daccu1_o1_c VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__a21oi_1
X_1682_ _0133_ _0611_ dsmod_daccu1_o1_c _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a31o_1
X_1683_ _0643_ _0612_ dsmod_daccu1_o0_c _0118_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and4b_1
X_1684_ _0133_ _0615_ dsmod_daccu1_o1_c _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a31o_1
X_1685_ dsmod_daccu1_o3_c _0635_ _0140_ _0612_ dsmod_daccu1_o2_c VGND VGND VPWR VPWR _0646_
+ sky130_fd_sc_hd__o2111a_1
X_1686_ _0147_ _0615_ dsmod_daccu1_o3_c _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a31o_1
X_1687_ _0636_ _0641_ _0645_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a31o_1
X_1688_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__inv_2
X_1689_ _0628_ _0634_ _0622_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or4_1
X_1690_ _0610_ _0613_ _0617_ _0626_ _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o2111a_1
X_1691_ dsmod_daccu1_o9_c _0607_ dsmod_daccu1_o9_c _0607_ VGND VGND VPWR VPWR _0652_
+ sky130_fd_sc_hd__o2bb2a_1
X_1692_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__inv_2
X_1693_ _0070_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__inv_2
X_1694_ dsmod_daccu1_o8_c VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__inv_2
X_1695_ _0579_ _0654_ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__o21a_1
X_1696_ _0585_ _0070_ dsmod_daccu1_o8_c _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a31o_1
X_1697_ _0653_ _0657_ _0606_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or3_1
X_1698_ dsmod_daccu1_o11_c _0601_ _0586_ _0136_ dsmod_daccu1_o10_c VGND VGND VPWR VPWR _0659_
+ sky130_fd_sc_hd__o2111a_1
X_1699_ dsmod_daccu1_o11_c _0601_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__a21oi_1
X_1700_ _0606_ _0609_ _0651_ _0658_ _0660_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__o221a_1
X_1701_ _0593_ _0594_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2_1
X_1702_ _0598_ _0599_ _0595_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or3_1
X_1703_ _0596_ _0600_ _0661_ _0662_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o311a_1
X_1704_ _0591_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__nor2_1
X_1705_ _0587_ _0154_ dsmod_daccu1_o14_c _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__a31o_1
X_1706_ _0584_ _0666_ net18 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a21o_1
X_1707_ _0575_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__clkbuf_4
X_1708_ net27 _0577_ _0583_ _0667_ _0668_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__o221a_1
X_1709_ _0815_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__clkbuf_4
X_1710_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__buf_2
X_1711_ _0584_ _0666_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nor2_1
X_1712_ _0576_ _0578_ _0667_ _0671_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o22a_1
X_1713_ _0670_ _0672_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__nor2_1
X_1714_ net18 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__clkbuf_2
X_1715_ _0591_ _0664_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and2_1
X_1716_ _0576_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_2
X_1717_ _0673_ _0665_ _0674_ _0675_ _0589_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o32a_1
X_1718_ _0670_ _0676_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nor2_1
X_1719_ _0675_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__buf_2
X_1720_ _0871_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__clkbuf_4
X_1721_ _0596_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__inv_2
X_1722_ _0598_ _0599_ _0661_ _0600_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o22a_1
X_1723_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__inv_2
X_1724_ net18 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__clkbuf_2
X_1725_ _0679_ _0680_ _0596_ _0681_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a221o_1
X_1726_ _0677_ dsmod_daccu1_o13_c _0678_ _0683_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__o211a_1
X_1727_ _0673_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__clkbuf_2
X_1728_ _0661_ _0600_ _0661_ _0600_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__a2bb2oi_1
X_1729_ _0577_ dsmod_daccu1_o12_c _0684_ _0685_ _0668_ VGND VGND VPWR VPWR _0206_
+ sky130_fd_sc_hd__o221a_1
X_1730_ _0653_ _0657_ _0651_ _0609_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o31a_1
X_1731_ _0605_ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor2_1
X_1732_ _0587_ _0136_ dsmod_daccu1_o10_c _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a31o_1
X_1733_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__inv_2
X_1734_ _0602_ _0689_ _0603_ _0688_ _0682_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__a221o_1
X_1735_ _0677_ dsmod_daccu1_o11_c _0678_ _0690_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__o211a_1
X_1736_ _0605_ _0686_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__and2_1
X_1737_ dsmod_daccu1_o10_c VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__inv_2
X_1738_ _0673_ _0687_ _0691_ _0675_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o32a_1
X_1739_ _0670_ _0693_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_1
X_1740_ _0579_ _0654_ _0655_ _0651_ _0657_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o32a_1
X_1741_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__inv_2
X_1742_ _0652_ _0694_ _0653_ _0695_ _0682_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a221o_1
X_1743_ _0677_ dsmod_daccu1_o9_c _0678_ _0696_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o211a_1
X_1744_ _0651_ _0657_ _0651_ _0657_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a2bb2oi_1
X_1745_ _0577_ dsmod_daccu1_o8_c _0684_ _0697_ _0668_ VGND VGND VPWR VPWR _0202_
+ sky130_fd_sc_hd__o221a_1
X_1746_ _0628_ _0634_ _0649_ _0625_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o31a_1
X_1747_ _0621_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__nor2_1
X_1748_ _0156_ _0616_ dsmod_daccu1_o6_c _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a31o_1
X_1749_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__inv_2
X_1750_ _0618_ _0701_ _0619_ _0700_ _0682_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__a221o_1
X_1751_ _0677_ dsmod_daccu1_o7_c _0872_ _0702_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__o211a_1
X_1752_ _0621_ _0698_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and2_1
X_1753_ dsmod_daccu1_o6_c VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__inv_2
X_1754_ _0673_ _0699_ _0703_ _0675_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o32a_1
X_1755_ _0670_ _0705_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__nor2_1
X_1756_ _0629_ _0631_ _0632_ _0649_ _0634_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o32a_1
X_1757_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__inv_2
X_1758_ _0627_ _0706_ _0628_ _0707_ _0682_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a221o_1
X_1759_ _0677_ dsmod_daccu1_o5_c _0872_ _0708_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__o211a_1
X_1760_ _0634_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__inv_2
X_1761_ _0649_ _0634_ _0648_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__o22a_1
X_1762_ _0871_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__clkbuf_4
X_1763_ _0577_ dsmod_daccu1_o4_c _0684_ _0710_ _0711_ VGND VGND VPWR VPWR _0198_
+ sky130_fd_sc_hd__o221a_1
X_1764_ _0645_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__inv_2
X_1765_ _0637_ _0631_ _0638_ _0712_ _0640_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__o32a_1
X_1766_ _0636_ _0713_ _0684_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a21oi_1
X_1767_ _0636_ _0713_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__o21ai_1
X_1768_ _0577_ dsmod_daccu1_o3_c _0872_ _0715_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__o211a_1
X_1769_ _0712_ _0640_ _0645_ _0641_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__o22a_1
X_1770_ _0675_ dsmod_daccu1_o2_c _0684_ _0716_ _0711_ VGND VGND VPWR VPWR _0196_
+ sky130_fd_sc_hd__o221a_1
X_1771_ _0118_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__inv_2
X_1772_ dsmod_daccu1_o0_c VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__inv_2
X_1773_ _0717_ _0631_ _0718_ _0643_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o31a_1
X_1774_ dsmod_daccu1_o1_c VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__inv_2
X_1775_ _0673_ _0644_ _0719_ _0576_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o32a_1
X_1776_ _0670_ _0721_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__nor2_1
X_1777_ _0717_ _0631_ net18 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or3_1
X_1778_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__inv_2
X_1779_ dsmod_daccu1_o0_c _0723_ _0718_ _0722_ _0711_ VGND VGND VPWR VPWR _0194_
+ sky130_fd_sc_hd__o221a_1
X_1780_ _0817_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__clkbuf_2
X_1781_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__clkinv_2
X_1782_ _0815_ _0795_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nor2_1
X_1783_ net28 _0725_ _0184_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__o21a_1
X_1784_ dsmod_dfetch__ctr_o0_c dsmod_dfetch__ctr_o1_c VGND VGND VPWR VPWR _0726_
+ sky130_fd_sc_hd__or2_1
X_1785_ dsmod_dfetch__ctr_o2_c _0726_ dsmod_dfetch__ctr_o3_c VGND VGND VPWR VPWR _0727_
+ sky130_fd_sc_hd__or3_1
X_1786_ dsmod_dfetch__ctr_o4_c _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__or2_1
X_1787_ dsmod_dfetch__ctr_o5_c _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__or2_1
X_1788_ dsmod_dfetch__ctr_o6_c _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__or2_1
X_1789_ fifo_dread__ptr_o3_c fifo_dwrite__ptr_o3_c _0010_ _0789_ VGND VGND VPWR VPWR _0731_
+ sky130_fd_sc_hd__o22a_1
X_1790_ fifo_dread__ptr_o1_c fifo_dwrite__ptr_o1_c _0008_ _0784_ VGND VGND VPWR VPWR _0732_
+ sky130_fd_sc_hd__o22a_1
X_1791_ _0731_ _0801_ _0800_ _0732_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__nor4_2
X_1792_ dsmod_dfetch__ctr_o7_c _0730_ net29 VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__or3_1
X_1793_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__clkbuf_2
X_1794_ _0734_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkinv_2
X_1795_ _0008_ _0799_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__or2_1
X_1796_ _0009_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__or2_1
X_1797_ fifo_dread__ptr_o3_c _0736_ fifo_dread__ptr_o3_c _0736_ VGND VGND VPWR VPWR _0020_
+ sky130_fd_sc_hd__o2bb2a_1
X_1798_ _0007_ _0020_ _0010_ _0734_ _0669_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a221oi_1
X_1799_ _0009_ _0735_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__a21bo_1
X_1800_ _0737_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_1801_ _0007_ _0012_ _0009_ _0734_ _0669_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a221oi_1
X_1802_ fifo_dread__ptr_o1_c fifo_dread__ptr_o0_c _0735_ VGND VGND VPWR VPWR _0013_
+ sky130_fd_sc_hd__o21ai_1
X_1803_ _0008_ _0734_ _0007_ _0013_ _0669_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__a221oi_1
X_1804_ fifo_dread__ptr_o0_c _0007_ _0799_ _0734_ _0563_ VGND VGND VPWR VPWR _0189_
+ sky130_fd_sc_hd__o221a_1
X_1805_ _0796_ _0724_ fifo_dwrite__ptr_o3_c _0725_ _0711_ VGND VGND VPWR VPWR _0188_
+ sky130_fd_sc_hd__o221a_1
X_1806_ _0793_ _0724_ fifo_dwrite__ptr_o2_c _0725_ _0711_ VGND VGND VPWR VPWR _0187_
+ sky130_fd_sc_hd__o221a_1
X_1807_ _0798_ _0724_ _0782_ _0725_ _0678_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__o221a_1
X_1808_ _0785_ _0724_ _0783_ _0725_ _0678_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__o221a_1
X_1809_ _0575_ _0006_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__and2_1
X_1810_ _0738_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_1811_ _0575_ _0005_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__and2_1
X_1812_ _0739_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_1813_ _0575_ _0004_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__and2_1
X_1814_ _0740_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
X_1815_ _0728_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__inv_2
X_1816_ dsmod_dfetch__ctr_o4_c _0727_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and2_1
X_1817_ _0741_ _0742_ _0668_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__o21a_1
X_1818_ _0727_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__inv_2
X_1819_ dsmod_dfetch__ctr_o2_c _0726_ dsmod_dfetch__ctr_o3_c VGND VGND VPWR VPWR _0744_
+ sky130_fd_sc_hd__o21a_1
X_1820_ _0743_ _0744_ _0668_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__o21a_1
X_1821_ _0815_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1822_ dsmod_dfetch__ctr_o2_c _0726_ dsmod_dfetch__ctr_o2_c _0726_ VGND VGND VPWR VPWR _0746_
+ sky130_fd_sc_hd__a2bb2oi_1
X_1823_ _0745_ _0746_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nor2_1
X_1824_ dsmod_dfetch__ctr_o0_c dsmod_dfetch__ctr_o1_c VGND VGND VPWR VPWR _0747_
+ sky130_fd_sc_hd__nand2_1
X_1825_ _0726_ _0747_ _0669_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__a21oi_1
X_1826_ _0745_ dsmod_dfetch__ctr_o0_c VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__nor2_1
X_1827_ fifo_dfifo__reg_o15_c_o15_c VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__inv_2
X_1828_ _0904_ _0492_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or2_4
X_1829_ _0870_ _0817_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a21oi_4
X_1830_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_2
X_1831_ _0749_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__clkbuf_2
X_1832_ _0748_ _0751_ _0908_ _0752_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__o22ai_1
X_1833_ fifo_dfifo__reg_o15_c_o14_c VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__inv_2
X_1834_ _0753_ _0751_ _0818_ _0752_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__o22ai_1
X_1835_ fifo_dfifo__reg_o15_c_o13_c VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__inv_2
X_1836_ _0754_ _0751_ _0821_ _0752_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__o22ai_1
X_1837_ fifo_dfifo__reg_o15_c_o12_c VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__inv_2
X_1838_ _0755_ _0751_ _0825_ _0752_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__o22ai_1
X_1839_ fifo_dfifo__reg_o15_c_o11_c VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__inv_2
X_1840_ _0756_ _0751_ _0829_ _0752_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__o22ai_1
X_1841_ fifo_dfifo__reg_o15_c_o10_c VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__inv_2
X_1842_ _0750_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__clkbuf_2
X_1843_ _0749_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__clkbuf_2
X_1844_ _0757_ _0758_ _0832_ _0759_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__o22ai_1
X_1845_ fifo_dfifo__reg_o15_c_o9_c VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__inv_2
X_1846_ _0760_ _0758_ _0837_ _0759_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o22ai_1
X_1847_ fifo_dfifo__reg_o15_c_o8_c VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__inv_2
X_1848_ _0761_ _0758_ _0840_ _0759_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o22ai_1
X_1849_ fifo_dfifo__reg_o15_c_o7_c VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__inv_2
X_1850_ _0762_ _0758_ _0844_ _0759_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__o22ai_1
X_1851_ fifo_dfifo__reg_o15_c_o6_c VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__inv_2
X_1852_ _0763_ _0758_ _0848_ _0759_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__o22ai_1
X_1853_ fifo_dfifo__reg_o15_c_o5_c VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__inv_2
X_1854_ _0750_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_2
X_1855_ _0749_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__clkbuf_2
X_1856_ _0764_ _0765_ _0851_ _0766_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__o22ai_1
X_1857_ fifo_dfifo__reg_o15_c_o4_c VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__inv_2
X_1858_ _0767_ _0765_ _0856_ _0766_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__o22ai_1
X_1859_ fifo_dfifo__reg_o15_c_o3_c VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__inv_2
X_1860_ _0768_ _0765_ _0859_ _0766_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__o22ai_1
X_1861_ fifo_dfifo__reg_o15_c_o2_c VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__inv_2
X_1862_ _0769_ _0765_ _0862_ _0766_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__o22ai_1
X_1863_ fifo_dfifo__reg_o15_c_o1_c VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__inv_2
X_1864_ _0770_ _0765_ _0865_ _0766_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o22ai_1
X_1865_ fifo_dfifo__reg_o15_c_o0_c VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__inv_2
X_1866_ _0771_ _0750_ _0868_ _0749_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__o22ai_1
X_1867_ _0745_ _0021_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__nor2_1
X_1868_ _0745_ _0022_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nor2_1
X_1869_ _0189_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__clkbuf_1
X_1870_ _0772_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
X_1871_ _0745_ _0023_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__nor2_1
X_1872_ dsmod_dfetch__ctr_o6_c _0729_ _0730_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a21bo_1
X_1873_ dsmod_dfetch__ctr_o7_c _0730_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__nor2_2
X_1874_ dsmod_dfetch__ctr_o7_c _0730_ _0011_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a21o_1
X_1875_ net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__inv_2
X_1876_ net19 net20 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__or2_1
X_1877_ _0773_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
X_1878_ dsmod_dfetch__ctr_o5_c _0728_ _0729_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a21bo_1
X_1879_ net19 net20 VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__and2_1
X_1880_ _0774_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
X_1881_ net20 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__clkbuf_1
X_1882_ _0775_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
X_1883_ net22 _0028_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__and2_1
X_1884_ _0776_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_1885_ net23 _0034_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__and2_1
X_1886_ _0777_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
X_1887_ _0581_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkinv_2
X_1888_ fifo_dfifo__reg_o9_c_o15_c VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__inv_2
X_1889_ _0778_ _0811_ _0810_ _0909_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o22ai_1
X_1890_ _0142_ _0144_ net24 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
X_1891_ _0157_ _0158_ net25 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
X_1892_ _0135_ _0137_ net24 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
X_1893_ _0154_ _0155_ net25 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
X_1894_ _0124_ _0128_ net24 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
X_1895_ _0151_ _0152_ net25 VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
X_1896_ _0069_ _0093_ net24 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_1
X_1897_ _0148_ _0149_ net25 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
X_1898_ _0127_ _0129_ net23 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
X_1899_ _0144_ _0145_ net24 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
X_1900_ _0143_ _0146_ net25 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
X_1901_ _0123_ _0126_ net23 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
X_1902_ _0141_ _0142_ net24 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
X_1903_ _0120_ _0122_ net23 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
X_1904_ _0092_ _0104_ net23 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_1
X_1905_ _0137_ _0138_ net24 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
X_1906_ _0136_ _0139_ net25 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
X_1907_ _0068_ _0081_ net23 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
X_1908_ _0134_ _0135_ net24 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_2
X_1909_ _0045_ _0057_ net23 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
X_1910_ _0103_ _0109_ net22 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_1
X_1911_ _0129_ _0130_ net23 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_1
X_1912_ _0128_ _0131_ net24 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
X_1913_ _0125_ _0132_ net25 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
X_1914_ _0091_ _0098_ net22 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
X_1915_ _0126_ _0127_ net23 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__mux2_1
X_1916_ _0080_ _0086_ net22 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_1
X_1917_ _0067_ _0075_ net22 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_1
X_1918_ _0121_ _0124_ net24 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
X_1919_ _0122_ _0123_ net23 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
X_1920_ _0056_ _0062_ net22 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
X_1921_ _0044_ _0051_ net22 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_1
X_1922_ _0119_ _0120_ net23 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
X_1923_ _0033_ _0039_ net22 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_1
X_1924_ _0109_ _0114_ net22 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_1
X_1925_ _0104_ _0115_ net23 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_1
X_1926_ _0093_ _0116_ net24 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
X_1927_ _0070_ _0117_ net25 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_1
X_1928_ _0098_ _0103_ net22 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
X_1929_ _0081_ _0092_ net23 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
X_1930_ _0086_ _0091_ net22 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
X_1931_ _0075_ _0080_ net22 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
X_1932_ _0046_ _0069_ net24 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_2
X_1933_ _0057_ _0068_ net23 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
X_1934_ _0062_ _0067_ net22 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
X_1935_ _0051_ _0056_ net22 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
X_1936_ _0034_ _0045_ net23 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_1
X_1937_ _0039_ _0044_ net22 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
X_1938_ _0028_ _0033_ net22 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
X_1939_ _0010_ _0020_ _0007_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_1
X_1940_ _0008_ _0013_ _0007_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_1
X_1941_ _0009_ _0012_ _0007_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_1
X_1942_ _0019_ _0016_ _0011_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_1
X_1943_ _0018_ _0017_ _0011_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_1
X_1944_ _0015_ _0014_ _0011_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
X_1945_ fifo_dfifo__reg_o0_c_o0_c fifo_dfifo__reg_o1_c_o0_c fifo_dfifo__reg_o2_c_o0_c
+ fifo_dfifo__reg_o3_c_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0110_
+ sky130_fd_sc_hd__mux4_1
X_1946_ fifo_dfifo__reg_o4_c_o0_c fifo_dfifo__reg_o5_c_o0_c fifo_dfifo__reg_o6_c_o0_c
+ fifo_dfifo__reg_o7_c_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0111_
+ sky130_fd_sc_hd__mux4_1
X_1947_ fifo_dfifo__reg_o8_c_o0_c fifo_dfifo__reg_o9_c_o0_c fifo_dfifo__reg_o10_c_o0_c
+ fifo_dfifo__reg_o11_c_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0112_
+ sky130_fd_sc_hd__mux4_1
X_1948_ fifo_dfifo__reg_o12_c_o0_c fifo_dfifo__reg_o13_c_o0_c fifo_dfifo__reg_o14_c_o0_c
+ fifo_dfifo__reg_o15_c_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0113_
+ sky130_fd_sc_hd__mux4_1
X_1949_ _0110_ _0111_ _0112_ _0113_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux4_2
X_1950_ fifo_dfifo__reg_o0_c_o1_c fifo_dfifo__reg_o1_c_o1_c fifo_dfifo__reg_o2_c_o1_c
+ fifo_dfifo__reg_o3_c_o1_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0105_
+ sky130_fd_sc_hd__mux4_1
X_1951_ fifo_dfifo__reg_o4_c_o1_c fifo_dfifo__reg_o5_c_o1_c fifo_dfifo__reg_o6_c_o1_c
+ fifo_dfifo__reg_o7_c_o1_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0106_
+ sky130_fd_sc_hd__mux4_2
X_1952_ fifo_dfifo__reg_o8_c_o1_c fifo_dfifo__reg_o9_c_o1_c fifo_dfifo__reg_o10_c_o1_c
+ fifo_dfifo__reg_o11_c_o1_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0107_
+ sky130_fd_sc_hd__mux4_1
X_1953_ fifo_dfifo__reg_o12_c_o1_c fifo_dfifo__reg_o13_c_o1_c fifo_dfifo__reg_o14_c_o1_c
+ fifo_dfifo__reg_o15_c_o1_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0108_
+ sky130_fd_sc_hd__mux4_1
X_1954_ _0105_ _0106_ _0107_ _0108_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux4_2
X_1955_ fifo_dfifo__reg_o0_c_o2_c fifo_dfifo__reg_o1_c_o2_c fifo_dfifo__reg_o2_c_o2_c
+ fifo_dfifo__reg_o3_c_o2_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0099_
+ sky130_fd_sc_hd__mux4_2
X_1956_ fifo_dfifo__reg_o4_c_o2_c fifo_dfifo__reg_o5_c_o2_c fifo_dfifo__reg_o6_c_o2_c
+ fifo_dfifo__reg_o7_c_o2_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0100_
+ sky130_fd_sc_hd__mux4_1
X_1957_ fifo_dfifo__reg_o8_c_o2_c fifo_dfifo__reg_o9_c_o2_c fifo_dfifo__reg_o10_c_o2_c
+ fifo_dfifo__reg_o11_c_o2_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0101_
+ sky130_fd_sc_hd__mux4_1
X_1958_ fifo_dfifo__reg_o12_c_o2_c fifo_dfifo__reg_o13_c_o2_c fifo_dfifo__reg_o14_c_o2_c
+ fifo_dfifo__reg_o15_c_o2_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0102_
+ sky130_fd_sc_hd__mux4_1
X_1959_ _0099_ _0100_ _0101_ _0102_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux4_2
X_1960_ fifo_dfifo__reg_o0_c_o3_c fifo_dfifo__reg_o1_c_o3_c fifo_dfifo__reg_o2_c_o3_c
+ fifo_dfifo__reg_o3_c_o3_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0094_
+ sky130_fd_sc_hd__mux4_2
X_1961_ fifo_dfifo__reg_o4_c_o3_c fifo_dfifo__reg_o5_c_o3_c fifo_dfifo__reg_o6_c_o3_c
+ fifo_dfifo__reg_o7_c_o3_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0095_
+ sky130_fd_sc_hd__mux4_1
X_1962_ fifo_dfifo__reg_o8_c_o3_c fifo_dfifo__reg_o9_c_o3_c fifo_dfifo__reg_o10_c_o3_c
+ fifo_dfifo__reg_o11_c_o3_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0096_
+ sky130_fd_sc_hd__mux4_1
X_1963_ fifo_dfifo__reg_o12_c_o3_c fifo_dfifo__reg_o13_c_o3_c fifo_dfifo__reg_o14_c_o3_c
+ fifo_dfifo__reg_o15_c_o3_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0097_
+ sky130_fd_sc_hd__mux4_1
X_1964_ _0094_ _0095_ _0096_ _0097_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux4_2
X_1965_ fifo_dfifo__reg_o0_c_o4_c fifo_dfifo__reg_o1_c_o4_c fifo_dfifo__reg_o2_c_o4_c
+ fifo_dfifo__reg_o3_c_o4_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0087_
+ sky130_fd_sc_hd__mux4_1
X_1966_ fifo_dfifo__reg_o4_c_o4_c fifo_dfifo__reg_o5_c_o4_c fifo_dfifo__reg_o6_c_o4_c
+ fifo_dfifo__reg_o7_c_o4_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0088_
+ sky130_fd_sc_hd__mux4_1
X_1967_ fifo_dfifo__reg_o8_c_o4_c fifo_dfifo__reg_o9_c_o4_c fifo_dfifo__reg_o10_c_o4_c
+ fifo_dfifo__reg_o11_c_o4_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0089_
+ sky130_fd_sc_hd__mux4_1
X_1968_ fifo_dfifo__reg_o12_c_o4_c fifo_dfifo__reg_o13_c_o4_c fifo_dfifo__reg_o14_c_o4_c
+ fifo_dfifo__reg_o15_c_o4_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0090_
+ sky130_fd_sc_hd__mux4_1
X_1969_ _0087_ _0088_ _0089_ _0090_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux4_2
X_1970_ fifo_dfifo__reg_o0_c_o5_c fifo_dfifo__reg_o1_c_o5_c fifo_dfifo__reg_o2_c_o5_c
+ fifo_dfifo__reg_o3_c_o5_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0082_
+ sky130_fd_sc_hd__mux4_2
X_1971_ fifo_dfifo__reg_o4_c_o5_c fifo_dfifo__reg_o5_c_o5_c fifo_dfifo__reg_o6_c_o5_c
+ fifo_dfifo__reg_o7_c_o5_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0083_
+ sky130_fd_sc_hd__mux4_1
X_1972_ fifo_dfifo__reg_o8_c_o5_c fifo_dfifo__reg_o9_c_o5_c fifo_dfifo__reg_o10_c_o5_c
+ fifo_dfifo__reg_o11_c_o5_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0084_
+ sky130_fd_sc_hd__mux4_1
X_1973_ fifo_dfifo__reg_o12_c_o5_c fifo_dfifo__reg_o13_c_o5_c fifo_dfifo__reg_o14_c_o5_c
+ fifo_dfifo__reg_o15_c_o5_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0085_
+ sky130_fd_sc_hd__mux4_1
X_1974_ _0082_ _0083_ _0084_ _0085_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux4_2
X_1975_ fifo_dfifo__reg_o0_c_o6_c fifo_dfifo__reg_o1_c_o6_c fifo_dfifo__reg_o2_c_o6_c
+ fifo_dfifo__reg_o3_c_o6_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0076_
+ sky130_fd_sc_hd__mux4_1
X_1976_ fifo_dfifo__reg_o4_c_o6_c fifo_dfifo__reg_o5_c_o6_c fifo_dfifo__reg_o6_c_o6_c
+ fifo_dfifo__reg_o7_c_o6_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0077_
+ sky130_fd_sc_hd__mux4_1
X_1977_ fifo_dfifo__reg_o8_c_o6_c fifo_dfifo__reg_o9_c_o6_c fifo_dfifo__reg_o10_c_o6_c
+ fifo_dfifo__reg_o11_c_o6_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0078_
+ sky130_fd_sc_hd__mux4_1
X_1978_ fifo_dfifo__reg_o12_c_o6_c fifo_dfifo__reg_o13_c_o6_c fifo_dfifo__reg_o14_c_o6_c
+ fifo_dfifo__reg_o15_c_o6_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0079_
+ sky130_fd_sc_hd__mux4_2
X_1979_ _0076_ _0077_ _0078_ _0079_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux4_1
X_1980_ fifo_dfifo__reg_o0_c_o7_c fifo_dfifo__reg_o1_c_o7_c fifo_dfifo__reg_o2_c_o7_c
+ fifo_dfifo__reg_o3_c_o7_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0071_
+ sky130_fd_sc_hd__mux4_1
X_1981_ fifo_dfifo__reg_o4_c_o7_c fifo_dfifo__reg_o5_c_o7_c fifo_dfifo__reg_o6_c_o7_c
+ fifo_dfifo__reg_o7_c_o7_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0072_
+ sky130_fd_sc_hd__mux4_1
X_1982_ fifo_dfifo__reg_o8_c_o7_c fifo_dfifo__reg_o9_c_o7_c fifo_dfifo__reg_o10_c_o7_c
+ fifo_dfifo__reg_o11_c_o7_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0073_
+ sky130_fd_sc_hd__mux4_1
X_1983_ fifo_dfifo__reg_o12_c_o7_c fifo_dfifo__reg_o13_c_o7_c fifo_dfifo__reg_o14_c_o7_c
+ fifo_dfifo__reg_o15_c_o7_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0074_
+ sky130_fd_sc_hd__mux4_1
X_1984_ _0071_ _0072_ _0073_ _0074_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__mux4_1
X_1985_ fifo_dfifo__reg_o0_c_o8_c fifo_dfifo__reg_o1_c_o8_c fifo_dfifo__reg_o2_c_o8_c
+ fifo_dfifo__reg_o3_c_o8_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0063_
+ sky130_fd_sc_hd__mux4_1
X_1986_ fifo_dfifo__reg_o4_c_o8_c fifo_dfifo__reg_o5_c_o8_c fifo_dfifo__reg_o6_c_o8_c
+ fifo_dfifo__reg_o7_c_o8_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0064_
+ sky130_fd_sc_hd__mux4_1
X_1987_ fifo_dfifo__reg_o8_c_o8_c fifo_dfifo__reg_o9_c_o8_c fifo_dfifo__reg_o10_c_o8_c
+ fifo_dfifo__reg_o11_c_o8_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0065_
+ sky130_fd_sc_hd__mux4_1
X_1988_ fifo_dfifo__reg_o12_c_o8_c fifo_dfifo__reg_o13_c_o8_c fifo_dfifo__reg_o14_c_o8_c
+ fifo_dfifo__reg_o15_c_o8_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0066_
+ sky130_fd_sc_hd__mux4_2
X_1989_ _0063_ _0064_ _0065_ _0066_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux4_1
X_1990_ fifo_dfifo__reg_o0_c_o9_c fifo_dfifo__reg_o1_c_o9_c fifo_dfifo__reg_o2_c_o9_c
+ fifo_dfifo__reg_o3_c_o9_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0058_
+ sky130_fd_sc_hd__mux4_1
X_1991_ fifo_dfifo__reg_o4_c_o9_c fifo_dfifo__reg_o5_c_o9_c fifo_dfifo__reg_o6_c_o9_c
+ fifo_dfifo__reg_o7_c_o9_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0059_
+ sky130_fd_sc_hd__mux4_1
X_1992_ fifo_dfifo__reg_o8_c_o9_c fifo_dfifo__reg_o9_c_o9_c fifo_dfifo__reg_o10_c_o9_c
+ fifo_dfifo__reg_o11_c_o9_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0060_
+ sky130_fd_sc_hd__mux4_1
X_1993_ fifo_dfifo__reg_o12_c_o9_c fifo_dfifo__reg_o13_c_o9_c fifo_dfifo__reg_o14_c_o9_c
+ fifo_dfifo__reg_o15_c_o9_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0061_
+ sky130_fd_sc_hd__mux4_1
X_1994_ _0058_ _0059_ _0060_ _0061_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux4_1
X_1995_ fifo_dfifo__reg_o0_c_o10_c fifo_dfifo__reg_o1_c_o10_c fifo_dfifo__reg_o2_c_o10_c
+ fifo_dfifo__reg_o3_c_o10_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0052_
+ sky130_fd_sc_hd__mux4_1
X_1996_ fifo_dfifo__reg_o4_c_o10_c fifo_dfifo__reg_o5_c_o10_c fifo_dfifo__reg_o6_c_o10_c
+ fifo_dfifo__reg_o7_c_o10_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0053_
+ sky130_fd_sc_hd__mux4_2
X_1997_ fifo_dfifo__reg_o8_c_o10_c fifo_dfifo__reg_o9_c_o10_c fifo_dfifo__reg_o10_c_o10_c
+ fifo_dfifo__reg_o11_c_o10_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0054_
+ sky130_fd_sc_hd__mux4_1
X_1998_ fifo_dfifo__reg_o12_c_o10_c fifo_dfifo__reg_o13_c_o10_c fifo_dfifo__reg_o14_c_o10_c
+ fifo_dfifo__reg_o15_c_o10_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0055_
+ sky130_fd_sc_hd__mux4_1
X_1999_ _0052_ _0053_ _0054_ _0055_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux4_1
X_2000_ fifo_dfifo__reg_o0_c_o11_c fifo_dfifo__reg_o1_c_o11_c fifo_dfifo__reg_o2_c_o11_c
+ fifo_dfifo__reg_o3_c_o11_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0047_
+ sky130_fd_sc_hd__mux4_1
X_2001_ fifo_dfifo__reg_o4_c_o11_c fifo_dfifo__reg_o5_c_o11_c fifo_dfifo__reg_o6_c_o11_c
+ fifo_dfifo__reg_o7_c_o11_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0048_
+ sky130_fd_sc_hd__mux4_1
X_2002_ fifo_dfifo__reg_o8_c_o11_c fifo_dfifo__reg_o9_c_o11_c fifo_dfifo__reg_o10_c_o11_c
+ fifo_dfifo__reg_o11_c_o11_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0049_
+ sky130_fd_sc_hd__mux4_1
X_2003_ fifo_dfifo__reg_o12_c_o11_c fifo_dfifo__reg_o13_c_o11_c fifo_dfifo__reg_o14_c_o11_c
+ fifo_dfifo__reg_o15_c_o11_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0050_
+ sky130_fd_sc_hd__mux4_1
X_2004_ _0047_ _0048_ _0049_ _0050_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux4_1
X_2005_ fifo_dfifo__reg_o0_c_o12_c fifo_dfifo__reg_o1_c_o12_c fifo_dfifo__reg_o2_c_o12_c
+ fifo_dfifo__reg_o3_c_o12_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0040_
+ sky130_fd_sc_hd__mux4_1
X_2006_ fifo_dfifo__reg_o4_c_o12_c fifo_dfifo__reg_o5_c_o12_c fifo_dfifo__reg_o6_c_o12_c
+ fifo_dfifo__reg_o7_c_o12_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0041_
+ sky130_fd_sc_hd__mux4_1
X_2007_ fifo_dfifo__reg_o8_c_o12_c fifo_dfifo__reg_o9_c_o12_c fifo_dfifo__reg_o10_c_o12_c
+ fifo_dfifo__reg_o11_c_o12_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0042_
+ sky130_fd_sc_hd__mux4_1
X_2008_ fifo_dfifo__reg_o12_c_o12_c fifo_dfifo__reg_o13_c_o12_c fifo_dfifo__reg_o14_c_o12_c
+ fifo_dfifo__reg_o15_c_o12_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0043_
+ sky130_fd_sc_hd__mux4_1
X_2009_ _0040_ _0041_ _0042_ _0043_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux4_1
X_2010_ fifo_dfifo__reg_o0_c_o13_c fifo_dfifo__reg_o1_c_o13_c fifo_dfifo__reg_o2_c_o13_c
+ fifo_dfifo__reg_o3_c_o13_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0035_
+ sky130_fd_sc_hd__mux4_1
X_2011_ fifo_dfifo__reg_o4_c_o13_c fifo_dfifo__reg_o5_c_o13_c fifo_dfifo__reg_o6_c_o13_c
+ fifo_dfifo__reg_o7_c_o13_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0036_
+ sky130_fd_sc_hd__mux4_1
X_2012_ fifo_dfifo__reg_o8_c_o13_c fifo_dfifo__reg_o9_c_o13_c fifo_dfifo__reg_o10_c_o13_c
+ fifo_dfifo__reg_o11_c_o13_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0037_
+ sky130_fd_sc_hd__mux4_1
X_2013_ fifo_dfifo__reg_o12_c_o13_c fifo_dfifo__reg_o13_c_o13_c fifo_dfifo__reg_o14_c_o13_c
+ fifo_dfifo__reg_o15_c_o13_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0038_
+ sky130_fd_sc_hd__mux4_1
X_2014_ _0035_ _0036_ _0037_ _0038_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux4_2
X_2015_ fifo_dfifo__reg_o0_c_o14_c fifo_dfifo__reg_o1_c_o14_c fifo_dfifo__reg_o2_c_o14_c
+ fifo_dfifo__reg_o3_c_o14_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0029_
+ sky130_fd_sc_hd__mux4_1
X_2016_ fifo_dfifo__reg_o4_c_o14_c fifo_dfifo__reg_o5_c_o14_c fifo_dfifo__reg_o6_c_o14_c
+ fifo_dfifo__reg_o7_c_o14_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0030_
+ sky130_fd_sc_hd__mux4_1
X_2017_ fifo_dfifo__reg_o8_c_o14_c fifo_dfifo__reg_o9_c_o14_c fifo_dfifo__reg_o10_c_o14_c
+ fifo_dfifo__reg_o11_c_o14_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0031_
+ sky130_fd_sc_hd__mux4_1
X_2018_ fifo_dfifo__reg_o12_c_o14_c fifo_dfifo__reg_o13_c_o14_c fifo_dfifo__reg_o14_c_o14_c
+ fifo_dfifo__reg_o15_c_o14_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0032_
+ sky130_fd_sc_hd__mux4_1
X_2019_ _0029_ _0030_ _0031_ _0032_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux4_2
X_2020_ fifo_dfifo__reg_o0_c_o15_c fifo_dfifo__reg_o1_c_o15_c fifo_dfifo__reg_o2_c_o15_c
+ fifo_dfifo__reg_o3_c_o15_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0024_
+ sky130_fd_sc_hd__mux4_1
X_2021_ fifo_dfifo__reg_o4_c_o15_c fifo_dfifo__reg_o5_c_o15_c fifo_dfifo__reg_o6_c_o15_c
+ fifo_dfifo__reg_o7_c_o15_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0025_
+ sky130_fd_sc_hd__mux4_1
X_2022_ fifo_dfifo__reg_o8_c_o15_c fifo_dfifo__reg_o9_c_o15_c fifo_dfifo__reg_o10_c_o15_c
+ fifo_dfifo__reg_o11_c_o15_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0026_
+ sky130_fd_sc_hd__mux4_1
X_2023_ fifo_dfifo__reg_o12_c_o15_c fifo_dfifo__reg_o13_c_o15_c fifo_dfifo__reg_o14_c_o15_c
+ fifo_dfifo__reg_o15_c_o15_c fifo_dfifo__reg_srdreg_o0_c_sq_o0_c fifo_dfifo__reg_srdreg_o0_c_sq_o1_c VGND VGND VPWR VPWR _0027_
+ sky130_fd_sc_hd__mux4_1
X_2024_ _0024_ _0025_ _0026_ _0027_ fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ fifo_dfifo__reg_srdreg_o0_c_sq_o3_c VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux4_1
X_2025_ clknet_leaf_29_clk_i _0000_ VGND VGND VPWR VPWR fifo_dfifo__reg_srdreg_o0_c_sq_o0_c
+ sky130_fd_sc_hd__dfxtp_4
X_2026_ clknet_leaf_30_clk_i _0001_ VGND VGND VPWR VPWR fifo_dfifo__reg_srdreg_o0_c_sq_o1_c
+ sky130_fd_sc_hd__dfxtp_4
X_2027_ clknet_leaf_29_clk_i _0002_ VGND VGND VPWR VPWR fifo_dfifo__reg_srdreg_o0_c_sq_o2_c
+ sky130_fd_sc_hd__dfxtp_4
X_2028_ clknet_leaf_29_clk_i _0003_ VGND VGND VPWR VPWR fifo_dfifo__reg_srdreg_o0_c_sq_o3_c
+ sky130_fd_sc_hd__dfxtp_4
X_2029_ clknet_leaf_1_clk_i _0160_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2030_ clknet_leaf_1_clk_i _0161_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2031_ clknet_leaf_5_clk_i _0162_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2032_ clknet_leaf_5_clk_i _0163_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2033_ clknet_leaf_5_clk_i _0164_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2034_ clknet_leaf_5_clk_i _0165_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2035_ clknet_leaf_9_clk_i _0166_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2036_ clknet_leaf_11_clk_i _0167_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2037_ clknet_leaf_11_clk_i _0168_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2038_ clknet_leaf_18_clk_i _0169_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2039_ clknet_leaf_18_clk_i _0170_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2040_ clknet_leaf_27_clk_i _0171_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2041_ clknet_leaf_28_clk_i _0172_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2042_ clknet_leaf_28_clk_i _0173_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2043_ clknet_leaf_28_clk_i _0174_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2044_ clknet_leaf_27_clk_i _0175_ VGND VGND VPWR VPWR fifo_dfifo__reg_o15_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2045_ clknet_leaf_29_clk_i _0176_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2046_ clknet_leaf_29_clk_i _0177_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2047_ clknet_leaf_29_clk_i _0178_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2048_ clknet_leaf_29_clk_i _0179_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2049_ clknet_leaf_30_clk_i _0180_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2050_ clknet_leaf_30_clk_i _0181_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2051_ clknet_leaf_30_clk_i _0182_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2052_ clknet_leaf_30_clk_i _0183_ VGND VGND VPWR VPWR dsmod_dfetch__ctr_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2053_ clknet_leaf_0_clk_i _0184_ VGND VGND VPWR VPWR fifo_dfifo__rdy__last
+ sky130_fd_sc_hd__dfxtp_1
X_2054_ clknet_leaf_0_clk_i _0185_ VGND VGND VPWR VPWR fifo_dwrite__ptr_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2055_ clknet_leaf_0_clk_i _0186_ VGND VGND VPWR VPWR fifo_dwrite__ptr_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2056_ clknet_leaf_0_clk_i _0187_ VGND VGND VPWR VPWR fifo_dwrite__ptr_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2057_ clknet_leaf_0_clk_i _0188_ VGND VGND VPWR VPWR fifo_dwrite__ptr_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2058_ clknet_leaf_29_clk_i _0189_ VGND VGND VPWR VPWR fifo_dread__ptr_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2059_ clknet_leaf_30_clk_i _0190_ VGND VGND VPWR VPWR fifo_dread__ptr_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2060_ clknet_leaf_30_clk_i _0191_ VGND VGND VPWR VPWR fifo_dread__ptr_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2061_ clknet_leaf_30_clk_i _0192_ VGND VGND VPWR VPWR fifo_dread__ptr_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2062_ clknet_leaf_30_clk_i _0193_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
X_2063_ clknet_leaf_20_clk_i _0194_ VGND VGND VPWR VPWR dsmod_daccu1_o0_c sky130_fd_sc_hd__dfxtp_1
X_2064_ clknet_leaf_20_clk_i _0195_ VGND VGND VPWR VPWR dsmod_daccu1_o1_c sky130_fd_sc_hd__dfxtp_1
X_2065_ clknet_leaf_16_clk_i _0196_ VGND VGND VPWR VPWR dsmod_daccu1_o2_c sky130_fd_sc_hd__dfxtp_1
X_2066_ clknet_leaf_16_clk_i _0197_ VGND VGND VPWR VPWR dsmod_daccu1_o3_c sky130_fd_sc_hd__dfxtp_1
X_2067_ clknet_leaf_20_clk_i _0198_ VGND VGND VPWR VPWR dsmod_daccu1_o4_c sky130_fd_sc_hd__dfxtp_1
X_2068_ clknet_leaf_20_clk_i _0199_ VGND VGND VPWR VPWR dsmod_daccu1_o5_c sky130_fd_sc_hd__dfxtp_1
X_2069_ clknet_leaf_21_clk_i _0200_ VGND VGND VPWR VPWR dsmod_daccu1_o6_c sky130_fd_sc_hd__dfxtp_1
X_2070_ clknet_leaf_20_clk_i _0201_ VGND VGND VPWR VPWR dsmod_daccu1_o7_c sky130_fd_sc_hd__dfxtp_1
X_2071_ clknet_leaf_22_clk_i _0202_ VGND VGND VPWR VPWR dsmod_daccu1_o8_c sky130_fd_sc_hd__dfxtp_1
X_2072_ clknet_leaf_21_clk_i _0203_ VGND VGND VPWR VPWR dsmod_daccu1_o9_c sky130_fd_sc_hd__dfxtp_1
X_2073_ clknet_leaf_21_clk_i _0204_ VGND VGND VPWR VPWR dsmod_daccu1_o10_c sky130_fd_sc_hd__dfxtp_1
X_2074_ clknet_leaf_22_clk_i _0205_ VGND VGND VPWR VPWR dsmod_daccu1_o11_c sky130_fd_sc_hd__dfxtp_1
X_2075_ clknet_leaf_22_clk_i _0206_ VGND VGND VPWR VPWR dsmod_daccu1_o12_c sky130_fd_sc_hd__dfxtp_1
X_2076_ clknet_leaf_22_clk_i _0207_ VGND VGND VPWR VPWR dsmod_daccu1_o13_c sky130_fd_sc_hd__dfxtp_1
X_2077_ clknet_leaf_22_clk_i _0208_ VGND VGND VPWR VPWR dsmod_daccu1_o14_c sky130_fd_sc_hd__dfxtp_1
X_2078_ clknet_leaf_21_clk_i _0209_ VGND VGND VPWR VPWR dsmod_daccu1_o15_c sky130_fd_sc_hd__dfxtp_1
X_2079_ clknet_leaf_21_clk_i _0210_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_2
X_2080_ clknet_leaf_1_clk_i _0211_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2081_ clknet_leaf_6_clk_i _0212_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2082_ clknet_leaf_7_clk_i _0213_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2083_ clknet_leaf_7_clk_i _0214_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2084_ clknet_leaf_7_clk_i _0215_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2085_ clknet_leaf_7_clk_i _0216_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2086_ clknet_leaf_12_clk_i _0217_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2087_ clknet_leaf_9_clk_i _0218_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2088_ clknet_leaf_12_clk_i _0219_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2089_ clknet_leaf_12_clk_i _0220_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2090_ clknet_leaf_11_clk_i _0221_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2091_ clknet_leaf_27_clk_i _0222_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2092_ clknet_leaf_28_clk_i _0223_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2093_ clknet_leaf_28_clk_i _0224_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2094_ clknet_leaf_28_clk_i _0225_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2095_ clknet_leaf_26_clk_i _0226_ VGND VGND VPWR VPWR fifo_dfifo__reg_o0_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2096_ clknet_leaf_2_clk_i _0227_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2097_ clknet_leaf_4_clk_i _0228_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2098_ clknet_leaf_4_clk_i _0229_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2099_ clknet_leaf_4_clk_i _0230_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2100_ clknet_leaf_4_clk_i _0231_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2101_ clknet_leaf_4_clk_i _0232_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2102_ clknet_leaf_13_clk_i _0233_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2103_ clknet_leaf_13_clk_i _0234_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2104_ clknet_leaf_12_clk_i _0235_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2105_ clknet_leaf_18_clk_i _0236_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2106_ clknet_leaf_18_clk_i _0237_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2107_ clknet_leaf_26_clk_i _0238_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2108_ clknet_leaf_27_clk_i _0239_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2109_ clknet_leaf_27_clk_i _0240_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2110_ clknet_leaf_28_clk_i _0241_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2111_ clknet_leaf_26_clk_i _0242_ VGND VGND VPWR VPWR fifo_dfifo__reg_o10_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2112_ clknet_leaf_2_clk_i _0243_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2113_ clknet_leaf_4_clk_i _0244_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2114_ clknet_leaf_4_clk_i _0245_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2115_ clknet_leaf_4_clk_i _0246_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2116_ clknet_leaf_6_clk_i _0247_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2117_ clknet_leaf_6_clk_i _0248_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2118_ clknet_leaf_13_clk_i _0249_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2119_ clknet_leaf_13_clk_i _0250_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2120_ clknet_leaf_12_clk_i _0251_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2121_ clknet_leaf_17_clk_i _0252_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2122_ clknet_leaf_18_clk_i _0253_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2123_ clknet_leaf_25_clk_i _0254_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2124_ clknet_leaf_25_clk_i _0255_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2125_ clknet_leaf_24_clk_i _0256_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2126_ clknet_leaf_24_clk_i _0257_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2127_ clknet_leaf_26_clk_i _0258_ VGND VGND VPWR VPWR fifo_dfifo__reg_o11_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2128_ clknet_leaf_1_clk_i _0259_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2129_ clknet_leaf_1_clk_i _0260_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2130_ clknet_leaf_5_clk_i _0261_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2131_ clknet_leaf_5_clk_i _0262_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2132_ clknet_leaf_5_clk_i _0263_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2133_ clknet_leaf_5_clk_i _0264_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2134_ clknet_leaf_10_clk_i _0265_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2135_ clknet_leaf_10_clk_i _0266_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2136_ clknet_leaf_3_clk_i _0267_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2137_ clknet_leaf_3_clk_i _0268_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2138_ clknet_leaf_3_clk_i _0269_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2139_ clknet_leaf_0_clk_i _0270_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2140_ clknet_leaf_29_clk_i _0271_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2141_ clknet_leaf_29_clk_i _0272_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2142_ clknet_leaf_29_clk_i _0273_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2143_ clknet_leaf_2_clk_i _0274_ VGND VGND VPWR VPWR fifo_dfifo__reg_o12_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2144_ clknet_leaf_1_clk_i _0275_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2145_ clknet_leaf_1_clk_i _0276_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2146_ clknet_leaf_5_clk_i _0277_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2147_ clknet_leaf_5_clk_i _0278_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2148_ clknet_leaf_5_clk_i _0279_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2149_ clknet_leaf_5_clk_i _0280_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2150_ clknet_leaf_10_clk_i _0281_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2151_ clknet_leaf_10_clk_i _0282_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2152_ clknet_leaf_10_clk_i _0283_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2153_ clknet_leaf_3_clk_i _0284_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2154_ clknet_leaf_3_clk_i _0285_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2155_ clknet_leaf_27_clk_i _0286_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2156_ clknet_leaf_29_clk_i _0287_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2157_ clknet_leaf_29_clk_i _0288_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2158_ clknet_leaf_29_clk_i _0289_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2159_ clknet_leaf_2_clk_i _0290_ VGND VGND VPWR VPWR fifo_dfifo__reg_o13_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2160_ clknet_leaf_2_clk_i _0291_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2161_ clknet_leaf_2_clk_i _0292_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2162_ clknet_leaf_4_clk_i _0293_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2163_ clknet_leaf_4_clk_i _0294_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2164_ clknet_leaf_4_clk_i _0295_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2165_ clknet_leaf_4_clk_i _0296_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2166_ clknet_leaf_10_clk_i _0297_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2167_ clknet_leaf_10_clk_i _0298_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2168_ clknet_leaf_10_clk_i _0299_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2169_ clknet_leaf_11_clk_i _0300_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2170_ clknet_leaf_3_clk_i _0301_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2171_ clknet_leaf_27_clk_i _0302_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2172_ clknet_leaf_27_clk_i _0303_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2173_ clknet_leaf_29_clk_i _0304_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2174_ clknet_leaf_29_clk_i _0305_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2175_ clknet_leaf_2_clk_i _0306_ VGND VGND VPWR VPWR fifo_dfifo__reg_o14_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2176_ clknet_leaf_1_clk_i _0307_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2177_ clknet_leaf_6_clk_i _0308_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2178_ clknet_leaf_7_clk_i _0309_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2179_ clknet_leaf_7_clk_i _0310_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2180_ clknet_leaf_7_clk_i _0311_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2181_ clknet_leaf_7_clk_i _0312_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2182_ clknet_leaf_12_clk_i _0313_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2183_ clknet_leaf_14_clk_i _0314_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2184_ clknet_leaf_12_clk_i _0315_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2185_ clknet_leaf_17_clk_i _0316_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2186_ clknet_leaf_12_clk_i _0317_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2187_ clknet_leaf_27_clk_i _0318_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2188_ clknet_leaf_28_clk_i _0319_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2189_ clknet_leaf_28_clk_i _0320_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2190_ clknet_leaf_28_clk_i _0321_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2191_ clknet_leaf_26_clk_i _0322_ VGND VGND VPWR VPWR fifo_dfifo__reg_o1_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2192_ clknet_leaf_2_clk_i _0323_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2193_ clknet_leaf_6_clk_i _0324_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2194_ clknet_leaf_7_clk_i _0325_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2195_ clknet_leaf_7_clk_i _0326_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2196_ clknet_leaf_6_clk_i _0327_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2197_ clknet_leaf_6_clk_i _0328_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2198_ clknet_leaf_12_clk_i _0329_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2199_ clknet_leaf_15_clk_i _0330_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2200_ clknet_leaf_12_clk_i _0331_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2201_ clknet_leaf_17_clk_i _0332_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2202_ clknet_leaf_12_clk_i _0333_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2203_ clknet_leaf_26_clk_i _0334_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2204_ clknet_leaf_25_clk_i _0335_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2205_ clknet_leaf_28_clk_i _0336_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2206_ clknet_leaf_28_clk_i _0337_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2207_ clknet_leaf_26_clk_i _0338_ VGND VGND VPWR VPWR fifo_dfifo__reg_o2_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2208_ clknet_leaf_2_clk_i _0339_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2209_ clknet_leaf_8_clk_i _0340_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2210_ clknet_leaf_7_clk_i _0341_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2211_ clknet_leaf_7_clk_i _0342_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2212_ clknet_leaf_8_clk_i _0343_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2213_ clknet_leaf_8_clk_i _0344_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2214_ clknet_leaf_13_clk_i _0345_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2215_ clknet_leaf_14_clk_i _0346_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2216_ clknet_leaf_13_clk_i _0347_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2217_ clknet_leaf_16_clk_i _0348_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2218_ clknet_leaf_15_clk_i _0349_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2219_ clknet_leaf_25_clk_i _0350_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2220_ clknet_leaf_24_clk_i _0351_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2221_ clknet_leaf_28_clk_i _0352_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2222_ clknet_leaf_24_clk_i _0353_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2223_ clknet_leaf_25_clk_i _0354_ VGND VGND VPWR VPWR fifo_dfifo__reg_o3_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2224_ clknet_leaf_3_clk_i _0355_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2225_ clknet_leaf_9_clk_i _0356_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2226_ clknet_leaf_8_clk_i _0357_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2227_ clknet_leaf_8_clk_i _0358_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2228_ clknet_leaf_9_clk_i _0359_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2229_ clknet_leaf_9_clk_i _0360_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2230_ clknet_leaf_14_clk_i _0361_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2231_ clknet_leaf_14_clk_i _0362_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2232_ clknet_leaf_15_clk_i _0363_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2233_ clknet_leaf_15_clk_i _0364_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2234_ clknet_leaf_15_clk_i _0365_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2235_ clknet_leaf_21_clk_i _0366_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2236_ clknet_leaf_23_clk_i _0367_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2237_ clknet_leaf_23_clk_i _0368_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2238_ clknet_leaf_23_clk_i _0369_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2239_ clknet_leaf_19_clk_i _0370_ VGND VGND VPWR VPWR fifo_dfifo__reg_o4_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2240_ clknet_leaf_26_clk_i _0371_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2241_ clknet_leaf_9_clk_i _0372_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2242_ clknet_leaf_8_clk_i _0373_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2243_ clknet_leaf_8_clk_i _0374_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2244_ clknet_leaf_8_clk_i _0375_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2245_ clknet_leaf_9_clk_i _0376_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2246_ clknet_leaf_14_clk_i _0377_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2247_ clknet_leaf_14_clk_i _0378_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2248_ clknet_leaf_15_clk_i _0379_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2249_ clknet_leaf_16_clk_i _0380_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2250_ clknet_leaf_15_clk_i _0381_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2251_ clknet_leaf_21_clk_i _0382_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2252_ clknet_leaf_23_clk_i _0383_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2253_ clknet_leaf_23_clk_i _0384_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2254_ clknet_leaf_23_clk_i _0385_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2255_ clknet_leaf_19_clk_i _0386_ VGND VGND VPWR VPWR fifo_dfifo__reg_o5_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2256_ clknet_leaf_2_clk_i _0387_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2257_ clknet_leaf_9_clk_i _0388_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2258_ clknet_leaf_9_clk_i _0389_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2259_ clknet_leaf_9_clk_i _0390_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2260_ clknet_leaf_9_clk_i _0391_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2261_ clknet_leaf_9_clk_i _0392_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2262_ clknet_leaf_15_clk_i _0393_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2263_ clknet_leaf_15_clk_i _0394_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2264_ clknet_leaf_15_clk_i _0395_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2265_ clknet_leaf_16_clk_i _0396_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2266_ clknet_leaf_17_clk_i _0397_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2267_ clknet_leaf_25_clk_i _0398_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2268_ clknet_leaf_23_clk_i _0399_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2269_ clknet_leaf_23_clk_i _0400_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2270_ clknet_leaf_23_clk_i _0401_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2271_ clknet_leaf_18_clk_i _0402_ VGND VGND VPWR VPWR fifo_dfifo__reg_o6_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2272_ clknet_leaf_26_clk_i _0403_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2273_ clknet_leaf_9_clk_i _0404_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2274_ clknet_leaf_8_clk_i _0405_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2275_ clknet_leaf_8_clk_i _0406_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2276_ clknet_leaf_9_clk_i _0407_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2277_ clknet_leaf_13_clk_i _0408_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2278_ clknet_leaf_14_clk_i _0409_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2279_ clknet_leaf_14_clk_i _0410_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2280_ clknet_leaf_15_clk_i _0411_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2281_ clknet_leaf_15_clk_i _0412_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2282_ clknet_leaf_15_clk_i _0413_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2283_ clknet_leaf_21_clk_i _0414_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2284_ clknet_leaf_23_clk_i _0415_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2285_ clknet_leaf_23_clk_i _0416_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2286_ clknet_leaf_23_clk_i _0417_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2287_ clknet_leaf_21_clk_i _0418_ VGND VGND VPWR VPWR fifo_dfifo__reg_o7_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2288_ clknet_leaf_2_clk_i _0419_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2289_ clknet_leaf_3_clk_i _0420_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2290_ clknet_leaf_3_clk_i _0421_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2291_ clknet_leaf_10_clk_i _0422_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2292_ clknet_leaf_10_clk_i _0423_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2293_ clknet_leaf_10_clk_i _0424_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2294_ clknet_leaf_11_clk_i _0425_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2295_ clknet_leaf_12_clk_i _0426_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2296_ clknet_leaf_12_clk_i _0427_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2297_ clknet_leaf_18_clk_i _0428_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2298_ clknet_leaf_18_clk_i _0429_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2299_ clknet_leaf_25_clk_i _0430_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2300_ clknet_leaf_25_clk_i _0431_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2301_ clknet_leaf_25_clk_i _0432_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2302_ clknet_leaf_25_clk_i _0433_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2303_ clknet_leaf_19_clk_i _0434_ VGND VGND VPWR VPWR fifo_dfifo__reg_o8_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
X_2304_ clknet_leaf_2_clk_i _0435_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o0_c
+ sky130_fd_sc_hd__dfxtp_1
X_2305_ clknet_leaf_8_clk_i _0436_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o1_c
+ sky130_fd_sc_hd__dfxtp_1
X_2306_ clknet_leaf_8_clk_i _0437_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o2_c
+ sky130_fd_sc_hd__dfxtp_1
X_2307_ clknet_leaf_8_clk_i _0438_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o3_c
+ sky130_fd_sc_hd__dfxtp_1
X_2308_ clknet_leaf_8_clk_i _0439_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o4_c
+ sky130_fd_sc_hd__dfxtp_1
X_2309_ clknet_leaf_13_clk_i _0440_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o5_c
+ sky130_fd_sc_hd__dfxtp_1
X_2310_ clknet_leaf_13_clk_i _0441_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o6_c
+ sky130_fd_sc_hd__dfxtp_1
X_2311_ clknet_leaf_13_clk_i _0442_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o7_c
+ sky130_fd_sc_hd__dfxtp_1
X_2312_ clknet_leaf_13_clk_i _0443_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o8_c
+ sky130_fd_sc_hd__dfxtp_1
X_2313_ clknet_leaf_18_clk_i _0444_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o9_c
+ sky130_fd_sc_hd__dfxtp_1
X_2314_ clknet_leaf_18_clk_i _0445_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o10_c
+ sky130_fd_sc_hd__dfxtp_1
X_2315_ clknet_leaf_25_clk_i _0446_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o11_c
+ sky130_fd_sc_hd__dfxtp_1
X_2316_ clknet_leaf_23_clk_i _0447_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o12_c
+ sky130_fd_sc_hd__dfxtp_1
X_2317_ clknet_leaf_24_clk_i _0448_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o13_c
+ sky130_fd_sc_hd__dfxtp_1
X_2318_ clknet_leaf_24_clk_i _0449_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o14_c
+ sky130_fd_sc_hd__dfxtp_1
X_2319_ clknet_leaf_26_clk_i _0450_ VGND VGND VPWR VPWR fifo_dfifo__reg_o9_c_o15_c
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_clk_i clk_i VGND VGND VPWR VPWR clknet_0_clk_i sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_0__f_clk_i clknet_0_clk_i VGND VGND VPWR VPWR clknet_2_0__leaf_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_1__f_clk_i clknet_0_clk_i VGND VGND VPWR VPWR clknet_2_1__leaf_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_2__f_clk_i clknet_0_clk_i VGND VGND VPWR VPWR clknet_2_2__leaf_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_3__f_clk_i clknet_0_clk_i VGND VGND VPWR VPWR clknet_2_3__leaf_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_0_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_0_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_10_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_10_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_11_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_11_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_12_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_12_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_13_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_13_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_14_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_15_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_15_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_16_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_16_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_17_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_17_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_18_clk_i clknet_2_3__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_18_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_19_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_19_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_1_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_1_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_20_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_20_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_21_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_21_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_22_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_22_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_23_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_23_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_24_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_24_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_25_clk_i clknet_2_2__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_25_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_26_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_27_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_27_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_28_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_29_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_29_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_2_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_2_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_30_clk_i clknet_2_0__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_30_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_3_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_3_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_4_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_4_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_5_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_5_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_6_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_6_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_7_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_7_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_8_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_8_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_9_clk_i clknet_2_1__leaf_clk_i VGND VGND VPWR VPWR clknet_leaf_9_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xinput1 fifo_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
Xinput10 fifo_i[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput11 fifo_i[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput12 fifo_i[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
Xinput13 fifo_i[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
Xinput14 fifo_i[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput15 fifo_i[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput16 fifo_i[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput17 fifo_rdy_i VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput18 mode_i VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput19 osr_i[0] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xinput2 fifo_i[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
Xinput20 osr_i[1] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput21 rst_n_i VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput22 volume_i[0] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_6
Xinput23 volume_i[1] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_6
Xinput24 volume_i[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_6
Xinput25 volume_i[3] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_6
Xinput3 fifo_i[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
Xinput4 fifo_i[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
Xinput5 fifo_i[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
Xinput6 fifo_i[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
Xinput7 fifo_i[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
Xinput8 fifo_i[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
Xinput9 fifo_i[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
Xoutput26 net26 VGND VGND VPWR VPWR ds_n_o sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR ds_o sky130_fd_sc_hd__buf_2
Xoutput28 net28 VGND VGND VPWR VPWR fifo_ack_o sky130_fd_sc_hd__buf_2
Xoutput29 net29 VGND VGND VPWR VPWR fifo_empty_o sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR fifo_full_o sky130_fd_sc_hd__buf_2
**.ends
.end
