** sch_path: /home/schippes/.xschem/xschem_library/xschem_sky130/xschem_verilog_import/spm.sch
**.subckt spm VGND VPWR clk p rst y
*+ x[31],x[30],x[29],x[28],x[27],x[26],x[25],x[24],x[23],x[22],x[21],x[20],x[19],x[18],x[17],x[16],x[15],x[14],x[13],x[12],x[11],x[10],x[9],x[8],x[7],x[6],x[5],x[4],x[3],x[2],x[1],x[0]
*.ipin VGND
*.ipin VPWR
*.ipin clk
*.opin p
*.ipin rst
*.ipin y
*.ipin
*+ x[31],x[30],x[29],x[28],x[27],x[26],x[25],x[24],x[23],x[22],x[21],x[20],x[19],x[18],x[17],x[16],x[15],x[14],x[13],x[12],x[11],x[10],x[9],x[8],x[7],x[6],x[5],x[4],x[3],x[2],x[1],x[0]
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_245_ net34 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__buf_2
X_246_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__dlymetal6s2s_1
X_247_ _098_ net2 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__and2_1
X_248_ csa0_dsc csa0_dy csa0_dsc csa0_dy VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__o2bb2a_1
X_249_ csa0_dsc csa0_dy _099_ _100_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a22o_1
X_250_ _099_ _100_ _099_ _100_ VGND VGND VPWR VPWR csa0_dhsum2 sky130_fd_sc_hd__o2bb2a_1
X_251_ _098_ net26 tcmp_dz VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__a21oi_1
X_252_ _098_ net26 tcmp_dz _101_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a31oi_1
X_253_ _101_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
X_254_ _098_ net13 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__and2_1
X_255_ genblk1_o1_c_dcsa_dsc genblk1_o1_c_dcsa_dy genblk1_o1_c_dcsa_dsc genblk1_o1_c_dcsa_dy VGND
+ VGND VPWR VPWR _103_ sky130_fd_sc_hd__o2bb2a_1
X_256_ genblk1_o1_c_dcsa_dsc genblk1_o1_c_dcsa_dy _102_ _103_ VGND VGND VPWR VPWR _011_
+ sky130_fd_sc_hd__a22o_1
X_257_ _102_ _103_ _102_ _103_ VGND VGND VPWR VPWR genblk1_o1_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_258_ _098_ net24 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__and2_1
X_259_ genblk1_o2_c_dcsa_dsc genblk1_o2_c_dcsa_dy genblk1_o2_c_dcsa_dsc genblk1_o2_c_dcsa_dy VGND
+ VGND VPWR VPWR _105_ sky130_fd_sc_hd__o2bb2a_1
X_260_ genblk1_o2_c_dcsa_dsc genblk1_o2_c_dcsa_dy _104_ _105_ VGND VGND VPWR VPWR _022_
+ sky130_fd_sc_hd__a22o_1
X_261_ _104_ _105_ _104_ _105_ VGND VGND VPWR VPWR genblk1_o2_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_262_ _097_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__clkbuf_1
X_263_ _106_ net27 VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__and2_1
X_264_ genblk1_o3_c_dcsa_dsc genblk1_o3_c_dcsa_dy genblk1_o3_c_dcsa_dsc genblk1_o3_c_dcsa_dy VGND
+ VGND VPWR VPWR _108_ sky130_fd_sc_hd__o2bb2a_1
X_265_ genblk1_o3_c_dcsa_dsc genblk1_o3_c_dcsa_dy _107_ _108_ VGND VGND VPWR VPWR _024_
+ sky130_fd_sc_hd__a22o_1
X_266_ _107_ _108_ _107_ _108_ VGND VGND VPWR VPWR genblk1_o3_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_267_ _106_ net28 VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__and2_1
X_268_ genblk1_o4_c_dcsa_dsc genblk1_o4_c_dcsa_dy genblk1_o4_c_dcsa_dsc genblk1_o4_c_dcsa_dy VGND
+ VGND VPWR VPWR _110_ sky130_fd_sc_hd__o2bb2a_1
X_269_ genblk1_o4_c_dcsa_dsc genblk1_o4_c_dcsa_dy _109_ _110_ VGND VGND VPWR VPWR _025_
+ sky130_fd_sc_hd__a22o_1
X_270_ _109_ _110_ _109_ _110_ VGND VGND VPWR VPWR genblk1_o4_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_271_ _106_ net29 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__and2_1
X_272_ genblk1_o5_c_dcsa_dsc genblk1_o5_c_dcsa_dy genblk1_o5_c_dcsa_dsc genblk1_o5_c_dcsa_dy VGND
+ VGND VPWR VPWR _112_ sky130_fd_sc_hd__o2bb2a_1
X_273_ genblk1_o5_c_dcsa_dsc genblk1_o5_c_dcsa_dy _111_ _112_ VGND VGND VPWR VPWR _026_
+ sky130_fd_sc_hd__a22o_1
X_274_ _111_ _112_ _111_ _112_ VGND VGND VPWR VPWR genblk1_o5_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_275_ _106_ net30 VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__and2_1
X_276_ genblk1_o6_c_dcsa_dsc genblk1_o6_c_dcsa_dy genblk1_o6_c_dcsa_dsc genblk1_o6_c_dcsa_dy VGND
+ VGND VPWR VPWR _114_ sky130_fd_sc_hd__o2bb2a_1
X_277_ genblk1_o6_c_dcsa_dsc genblk1_o6_c_dcsa_dy _113_ _114_ VGND VGND VPWR VPWR _027_
+ sky130_fd_sc_hd__a22o_1
X_278_ _113_ _114_ _113_ _114_ VGND VGND VPWR VPWR genblk1_o6_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_279_ _106_ net31 VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and2_1
X_280_ genblk1_o7_c_dcsa_dsc genblk1_o7_c_dcsa_dy genblk1_o7_c_dcsa_dsc genblk1_o7_c_dcsa_dy VGND
+ VGND VPWR VPWR _116_ sky130_fd_sc_hd__o2bb2a_1
X_281_ genblk1_o7_c_dcsa_dsc genblk1_o7_c_dcsa_dy _115_ _116_ VGND VGND VPWR VPWR _028_
+ sky130_fd_sc_hd__a22o_1
X_282_ _115_ _116_ _115_ _116_ VGND VGND VPWR VPWR genblk1_o7_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_283_ net34 VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__clkbuf_1
X_284_ _117_ net32 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__and2_1
X_285_ genblk1_o8_c_dcsa_dsc genblk1_o8_c_dcsa_dy genblk1_o8_c_dcsa_dsc genblk1_o8_c_dcsa_dy VGND
+ VGND VPWR VPWR _119_ sky130_fd_sc_hd__o2bb2a_1
X_286_ genblk1_o8_c_dcsa_dsc genblk1_o8_c_dcsa_dy _118_ _119_ VGND VGND VPWR VPWR _029_
+ sky130_fd_sc_hd__a22o_1
X_287_ _118_ _119_ _118_ _119_ VGND VGND VPWR VPWR genblk1_o8_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_288_ _117_ net33 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__and2_1
X_289_ genblk1_o9_c_dcsa_dsc genblk1_o10_c_dcsa_dsum genblk1_o9_c_dcsa_dsc genblk1_o10_c_dcsa_dsum
+ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__o2bb2a_1
X_290_ genblk1_o9_c_dcsa_dsc genblk1_o10_c_dcsa_dsum _120_ _121_ VGND VGND VPWR VPWR _030_
+ sky130_fd_sc_hd__a22o_1
X_291_ _120_ _121_ _120_ _121_ VGND VGND VPWR VPWR genblk1_o9_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_292_ _117_ net3 VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__and2_1
X_293_ genblk1_o10_c_dcsa_dsc genblk1_o10_c_dcsa_dy genblk1_o10_c_dcsa_dsc genblk1_o10_c_dcsa_dy
+ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__o2bb2a_1
X_294_ genblk1_o10_c_dcsa_dsc genblk1_o10_c_dcsa_dy _122_ _123_ VGND VGND VPWR VPWR _001_
+ sky130_fd_sc_hd__a22o_1
X_295_ _122_ _123_ _122_ _123_ VGND VGND VPWR VPWR genblk1_o10_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_296_ _117_ net4 VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__and2_1
X_297_ genblk1_o11_c_dcsa_dsc genblk1_o11_c_dcsa_dy genblk1_o11_c_dcsa_dsc genblk1_o11_c_dcsa_dy
+ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__o2bb2a_1
X_298_ genblk1_o11_c_dcsa_dsc genblk1_o11_c_dcsa_dy _124_ _125_ VGND VGND VPWR VPWR _002_
+ sky130_fd_sc_hd__a22o_1
X_299_ _124_ _125_ _124_ _125_ VGND VGND VPWR VPWR genblk1_o11_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_300_ _117_ net5 VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__and2_1
X_301_ genblk1_o12_c_dcsa_dsc genblk1_o12_c_dcsa_dy genblk1_o12_c_dcsa_dsc genblk1_o12_c_dcsa_dy
+ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__o2bb2a_1
X_302_ genblk1_o12_c_dcsa_dsc genblk1_o12_c_dcsa_dy _126_ _127_ VGND VGND VPWR VPWR _003_
+ sky130_fd_sc_hd__a22o_1
X_303_ _126_ _127_ _126_ _127_ VGND VGND VPWR VPWR genblk1_o12_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_304_ net34 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__clkbuf_1
X_305_ _128_ net6 VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__and2_1
X_306_ genblk1_o13_c_dcsa_dsc genblk1_o13_c_dcsa_dy genblk1_o13_c_dcsa_dsc genblk1_o13_c_dcsa_dy
+ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__o2bb2a_1
X_307_ genblk1_o13_c_dcsa_dsc genblk1_o13_c_dcsa_dy _129_ _130_ VGND VGND VPWR VPWR _004_
+ sky130_fd_sc_hd__a22o_1
X_308_ _129_ _130_ _129_ _130_ VGND VGND VPWR VPWR genblk1_o13_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_309_ _128_ net7 VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and2_1
X_310_ genblk1_o14_c_dcsa_dsc genblk1_o14_c_dcsa_dy genblk1_o14_c_dcsa_dsc genblk1_o14_c_dcsa_dy
+ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o2bb2a_1
X_311_ genblk1_o14_c_dcsa_dsc genblk1_o14_c_dcsa_dy _131_ _132_ VGND VGND VPWR VPWR _005_
+ sky130_fd_sc_hd__a22o_1
X_312_ _131_ _132_ _131_ _132_ VGND VGND VPWR VPWR genblk1_o14_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_313_ _128_ net8 VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__and2_1
X_314_ genblk1_o15_c_dcsa_dsc genblk1_o15_c_dcsa_dy genblk1_o15_c_dcsa_dsc genblk1_o15_c_dcsa_dy
+ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__o2bb2a_1
X_315_ genblk1_o15_c_dcsa_dsc genblk1_o15_c_dcsa_dy _133_ _134_ VGND VGND VPWR VPWR _006_
+ sky130_fd_sc_hd__a22o_1
X_316_ _133_ _134_ _133_ _134_ VGND VGND VPWR VPWR genblk1_o15_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_317_ _128_ net9 VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and2_1
X_318_ genblk1_o16_c_dcsa_dsc genblk1_o16_c_dcsa_dy genblk1_o16_c_dcsa_dsc genblk1_o16_c_dcsa_dy
+ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__o2bb2a_1
X_319_ genblk1_o16_c_dcsa_dsc genblk1_o16_c_dcsa_dy _135_ _136_ VGND VGND VPWR VPWR _007_
+ sky130_fd_sc_hd__a22o_1
X_320_ _135_ _136_ _135_ _136_ VGND VGND VPWR VPWR genblk1_o16_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_321_ _128_ net10 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__and2_1
X_322_ genblk1_o17_c_dcsa_dsc genblk1_o17_c_dcsa_dy genblk1_o17_c_dcsa_dsc genblk1_o17_c_dcsa_dy
+ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__o2bb2a_1
X_323_ genblk1_o17_c_dcsa_dsc genblk1_o17_c_dcsa_dy _137_ _138_ VGND VGND VPWR VPWR _008_
+ sky130_fd_sc_hd__a22o_1
X_324_ _137_ _138_ _137_ _138_ VGND VGND VPWR VPWR genblk1_o17_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_325_ net34 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__clkbuf_1
X_326_ _139_ net11 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__and2_1
X_327_ genblk1_o18_c_dcsa_dsc genblk1_o18_c_dcsa_dy genblk1_o18_c_dcsa_dsc genblk1_o18_c_dcsa_dy
+ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__o2bb2a_1
X_328_ genblk1_o18_c_dcsa_dsc genblk1_o18_c_dcsa_dy _140_ _141_ VGND VGND VPWR VPWR _009_
+ sky130_fd_sc_hd__a22o_1
X_329_ _140_ _141_ _140_ _141_ VGND VGND VPWR VPWR genblk1_o18_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_330_ _139_ net12 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__and2_1
X_331_ genblk1_o19_c_dcsa_dsc genblk1_o19_c_dcsa_dy genblk1_o19_c_dcsa_dsc genblk1_o19_c_dcsa_dy
+ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__o2bb2a_1
X_332_ genblk1_o19_c_dcsa_dsc genblk1_o19_c_dcsa_dy _142_ _143_ VGND VGND VPWR VPWR _010_
+ sky130_fd_sc_hd__a22o_1
X_333_ _142_ _143_ _142_ _143_ VGND VGND VPWR VPWR genblk1_o19_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_334_ _139_ net14 VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__and2_1
X_335_ genblk1_o20_c_dcsa_dsc genblk1_o20_c_dcsa_dy genblk1_o20_c_dcsa_dsc genblk1_o20_c_dcsa_dy
+ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__o2bb2a_1
X_336_ genblk1_o20_c_dcsa_dsc genblk1_o20_c_dcsa_dy _144_ _145_ VGND VGND VPWR VPWR _012_
+ sky130_fd_sc_hd__a22o_1
X_337_ _144_ _145_ _144_ _145_ VGND VGND VPWR VPWR genblk1_o20_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_338_ _139_ net15 VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__and2_1
X_339_ genblk1_o21_c_dcsa_dsc genblk1_o21_c_dcsa_dy genblk1_o21_c_dcsa_dsc genblk1_o21_c_dcsa_dy
+ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__o2bb2a_1
X_340_ genblk1_o21_c_dcsa_dsc genblk1_o21_c_dcsa_dy _146_ _147_ VGND VGND VPWR VPWR _013_
+ sky130_fd_sc_hd__a22o_1
X_341_ _146_ _147_ _146_ _147_ VGND VGND VPWR VPWR genblk1_o21_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_342_ _139_ net16 VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and2_1
X_343_ genblk1_o22_c_dcsa_dsc genblk1_o22_c_dcsa_dy genblk1_o22_c_dcsa_dsc genblk1_o22_c_dcsa_dy
+ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__o2bb2a_1
X_344_ genblk1_o22_c_dcsa_dsc genblk1_o22_c_dcsa_dy _148_ _149_ VGND VGND VPWR VPWR _014_
+ sky130_fd_sc_hd__a22o_1
X_345_ _148_ _149_ _148_ _149_ VGND VGND VPWR VPWR genblk1_o22_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_346_ net34 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__clkbuf_1
X_347_ _150_ net17 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__and2_1
X_348_ genblk1_o23_c_dcsa_dsc genblk1_o23_c_dcsa_dy genblk1_o23_c_dcsa_dsc genblk1_o23_c_dcsa_dy
+ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__o2bb2a_1
X_349_ genblk1_o23_c_dcsa_dsc genblk1_o23_c_dcsa_dy _151_ _152_ VGND VGND VPWR VPWR _015_
+ sky130_fd_sc_hd__a22o_1
X_350_ _151_ _152_ _151_ _152_ VGND VGND VPWR VPWR genblk1_o23_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_351_ _150_ net18 VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and2_1
X_352_ genblk1_o24_c_dcsa_dsc genblk1_o24_c_dcsa_dy genblk1_o24_c_dcsa_dsc genblk1_o24_c_dcsa_dy
+ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__o2bb2a_1
X_353_ genblk1_o24_c_dcsa_dsc genblk1_o24_c_dcsa_dy _153_ _154_ VGND VGND VPWR VPWR _016_
+ sky130_fd_sc_hd__a22o_1
X_354_ _153_ _154_ _153_ _154_ VGND VGND VPWR VPWR genblk1_o24_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_355_ _150_ net19 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__and2_1
X_356_ genblk1_o25_c_dcsa_dsc genblk1_o25_c_dcsa_dy genblk1_o25_c_dcsa_dsc genblk1_o25_c_dcsa_dy
+ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__o2bb2a_1
X_357_ genblk1_o25_c_dcsa_dsc genblk1_o25_c_dcsa_dy _155_ _156_ VGND VGND VPWR VPWR _017_
+ sky130_fd_sc_hd__a22o_1
X_358_ _155_ _156_ _155_ _156_ VGND VGND VPWR VPWR genblk1_o25_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_359_ _150_ net20 VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__and2_1
X_360_ genblk1_o26_c_dcsa_dsc genblk1_o26_c_dcsa_dy genblk1_o26_c_dcsa_dsc genblk1_o26_c_dcsa_dy
+ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__o2bb2a_1
X_361_ genblk1_o26_c_dcsa_dsc genblk1_o26_c_dcsa_dy _157_ _158_ VGND VGND VPWR VPWR _018_
+ sky130_fd_sc_hd__a22o_1
X_362_ _157_ _158_ _157_ _158_ VGND VGND VPWR VPWR genblk1_o26_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_363_ _150_ net21 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__and2_1
X_364_ genblk1_o27_c_dcsa_dsc genblk1_o27_c_dcsa_dy genblk1_o27_c_dcsa_dsc genblk1_o27_c_dcsa_dy
+ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__o2bb2a_1
X_365_ genblk1_o27_c_dcsa_dsc genblk1_o27_c_dcsa_dy _159_ _160_ VGND VGND VPWR VPWR _019_
+ sky130_fd_sc_hd__a22o_1
X_366_ _159_ _160_ _159_ _160_ VGND VGND VPWR VPWR genblk1_o27_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_367_ _097_ net22 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__and2_1
X_368_ genblk1_o28_c_dcsa_dsc genblk1_o28_c_dcsa_dy genblk1_o28_c_dcsa_dsc genblk1_o28_c_dcsa_dy
+ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__o2bb2a_1
X_369_ genblk1_o28_c_dcsa_dsc genblk1_o28_c_dcsa_dy _161_ _162_ VGND VGND VPWR VPWR _020_
+ sky130_fd_sc_hd__a22o_1
X_370_ _161_ _162_ _161_ _162_ VGND VGND VPWR VPWR genblk1_o28_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_371_ _097_ net23 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__and2_1
X_372_ genblk1_o29_c_dcsa_dsc genblk1_o29_c_dcsa_dy genblk1_o29_c_dcsa_dsc genblk1_o29_c_dcsa_dy
+ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__o2bb2a_1
X_373_ genblk1_o29_c_dcsa_dsc genblk1_o29_c_dcsa_dy _163_ _164_ VGND VGND VPWR VPWR _021_
+ sky130_fd_sc_hd__a22o_1
X_374_ _163_ _164_ _163_ _164_ VGND VGND VPWR VPWR genblk1_o29_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_375_ _097_ net25 VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__and2_1
X_376_ genblk1_o30_c_dcsa_dsc genblk1_o30_c_dcsa_dy genblk1_o30_c_dcsa_dsc genblk1_o30_c_dcsa_dy
+ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__o2bb2a_1
X_377_ genblk1_o30_c_dcsa_dsc genblk1_o30_c_dcsa_dy _165_ _166_ VGND VGND VPWR VPWR _023_
+ sky130_fd_sc_hd__a22o_1
X_378_ _165_ _166_ _165_ _166_ VGND VGND VPWR VPWR genblk1_o30_c_dcsa_dhsum2
+ sky130_fd_sc_hd__o2bb2a_1
X_379_ net1 VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__inv_2
X_380_ _167_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_2
X_381_ _033_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__clkbuf_1
X_382_ _168_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__clkbuf_1
X_383_ _033_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__clkbuf_1
X_384_ _169_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
X_385_ _033_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__clkbuf_1
X_386_ _170_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__clkbuf_1
X_387_ _033_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__clkbuf_1
X_388_ _171_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__clkbuf_1
X_389_ _167_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__dlymetal6s2s_1
X_390_ _172_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__dlymetal6s2s_1
X_391_ _173_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__clkbuf_1
X_392_ _174_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__clkbuf_1
X_393_ _173_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__clkbuf_1
X_394_ _175_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__clkbuf_1
X_395_ _173_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__clkbuf_1
X_396_ _176_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__clkbuf_1
X_397_ _173_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__clkbuf_1
X_398_ _177_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__clkbuf_1
X_399_ _173_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__clkbuf_1
X_400_ _178_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__clkbuf_1
X_401_ _167_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__dlymetal6s2s_1
X_402_ _179_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__dlymetal6s2s_1
X_403_ _180_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__clkbuf_1
X_404_ _181_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__clkbuf_1
X_405_ _180_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__clkbuf_1
X_406_ _182_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__clkbuf_1
X_407_ _180_ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__clkbuf_1
X_408_ _183_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__clkbuf_1
X_409_ _180_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__clkbuf_1
X_410_ _184_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__clkbuf_1
X_411_ _180_ VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__clkbuf_1
X_412_ _185_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__clkbuf_1
X_413_ _179_ VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__dlymetal6s2s_1
X_414_ _186_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__clkbuf_1
X_415_ _187_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__clkbuf_1
X_416_ _186_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__clkbuf_1
X_417_ _188_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__clkbuf_1
X_418_ _186_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__clkbuf_1
X_419_ _189_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__clkbuf_1
X_420_ _186_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__clkbuf_1
X_421_ _190_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkbuf_1
X_422_ _186_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__clkbuf_1
X_423_ _191_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__clkbuf_1
X_424_ _179_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__clkbuf_2
X_425_ _192_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__clkbuf_1
X_426_ _193_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__clkbuf_1
X_427_ _192_ VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__clkbuf_1
X_428_ _194_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__clkbuf_1
X_429_ _192_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__clkbuf_1
X_430_ _195_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__clkbuf_1
X_431_ _192_ VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__clkbuf_1
X_432_ _196_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__clkbuf_1
X_433_ _192_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__clkbuf_1
X_434_ _197_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__clkbuf_1
X_435_ _179_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__dlymetal6s2s_1
X_436_ _198_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__clkbuf_1
X_437_ _199_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__clkbuf_1
X_438_ _198_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__clkbuf_1
X_439_ _200_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__clkbuf_1
X_440_ _198_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__clkbuf_1
X_441_ _201_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__clkbuf_1
X_442_ _198_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__clkbuf_1
X_443_ _202_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__clkbuf_1
X_444_ _198_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__clkbuf_1
X_445_ _203_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__clkbuf_1
X_446_ _179_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__dlymetal6s2s_1
X_447_ _204_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__clkbuf_1
X_448_ _205_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__clkbuf_1
X_449_ _204_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__clkbuf_1
X_450_ _206_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__clkbuf_1
X_451_ _204_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__clkbuf_1
X_452_ _207_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__clkbuf_1
X_453_ _204_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__clkbuf_1
X_454_ _208_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__clkbuf_1
X_455_ _204_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__clkbuf_1
X_456_ _209_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__clkbuf_1
X_457_ _167_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__clkbuf_2
X_458_ _210_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__dlymetal6s2s_1
X_459_ _211_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__clkbuf_1
X_460_ _212_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__clkbuf_1
X_461_ _211_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__clkbuf_1
X_462_ _213_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__clkbuf_1
X_463_ _211_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__clkbuf_1
X_464_ _214_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__clkbuf_1
X_465_ _211_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__clkbuf_1
X_466_ _215_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__clkbuf_1
X_467_ _211_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__clkbuf_1
X_468_ _216_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__clkbuf_1
X_469_ _210_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__dlymetal6s2s_1
X_470_ _217_ VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__clkbuf_1
X_471_ _218_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__clkbuf_1
X_472_ _217_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__clkbuf_1
X_473_ _219_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__clkbuf_1
X_474_ _217_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__clkbuf_1
X_475_ _220_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__clkbuf_1
X_476_ _217_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__clkbuf_1
X_477_ _221_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__clkbuf_1
X_478_ _217_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__clkbuf_1
X_479_ _222_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__clkbuf_1
X_480_ _210_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__clkbuf_2
X_481_ _223_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__clkbuf_1
X_482_ _224_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__clkbuf_1
X_483_ _223_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__clkbuf_1
X_484_ _225_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__clkbuf_1
X_485_ _223_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__clkbuf_1
X_486_ _226_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__clkbuf_1
X_487_ _223_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__clkbuf_1
X_488_ _227_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__clkbuf_1
X_489_ _223_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__clkbuf_1
X_490_ _228_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__clkbuf_1
X_491_ _210_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__dlymetal6s2s_1
X_492_ _229_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__clkbuf_1
X_493_ _230_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__clkbuf_1
X_494_ _229_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__clkbuf_1
X_495_ _231_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__clkbuf_1
X_496_ _229_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__clkbuf_1
X_497_ _232_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__clkbuf_1
X_498_ _229_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__clkbuf_1
X_499_ _233_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__clkbuf_1
X_500_ _229_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__clkbuf_1
X_501_ _234_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__clkbuf_1
X_502_ _210_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__dlymetal6s2s_1
X_503_ _235_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__clkbuf_1
X_504_ _236_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__clkbuf_1
X_505_ _235_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__clkbuf_1
X_506_ _237_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__clkbuf_1
X_507_ _235_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__clkbuf_1
X_508_ _238_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__clkbuf_1
X_509_ _235_ VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__clkbuf_1
X_510_ _239_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__clkbuf_1
X_511_ _235_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__clkbuf_1
X_512_ _240_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__clkbuf_1
X_513_ _172_ VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__clkbuf_1
X_514_ _241_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__clkbuf_1
X_515_ _172_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__clkbuf_1
X_516_ _242_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__clkbuf_1
X_517_ _172_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__clkbuf_1
X_518_ _243_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__clkbuf_1
X_519_ _172_ VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__clkbuf_1
X_520_ _244_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__clkbuf_1
X_521_ clknet_3_0_0_clk _000_ _033_ VGND VGND VPWR VPWR csa0_dsc sky130_fd_sc_hd__dfrtp_1
X_522_ clknet_3_0_0_clk csa0_dhsum2 _034_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfrtp_1
X_523_ clknet_3_1_0_clk _032_ _035_ VGND VGND VPWR VPWR tcmp_dz sky130_fd_sc_hd__dfrtp_1
X_524_ clknet_3_1_0_clk _031_ _036_ VGND VGND VPWR VPWR genblk1_o30_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_525_ clknet_3_0_0_clk _011_ _037_ VGND VGND VPWR VPWR genblk1_o1_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_526_ clknet_3_0_0_clk genblk1_o1_c_dcsa_dhsum2 _038_ VGND VGND VPWR VPWR csa0_dy
+ sky130_fd_sc_hd__dfrtp_1
X_527_ clknet_3_0_0_clk _022_ _039_ VGND VGND VPWR VPWR genblk1_o2_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_528_ clknet_3_0_0_clk genblk1_o2_c_dcsa_dhsum2 _040_ VGND VGND VPWR VPWR genblk1_o1_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_529_ clknet_3_0_0_clk _024_ _041_ VGND VGND VPWR VPWR genblk1_o3_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_530_ clknet_3_0_0_clk genblk1_o3_c_dcsa_dhsum2 _042_ VGND VGND VPWR VPWR genblk1_o2_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_531_ clknet_3_2_0_clk _025_ _043_ VGND VGND VPWR VPWR genblk1_o4_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_532_ clknet_3_0_0_clk genblk1_o4_c_dcsa_dhsum2 _044_ VGND VGND VPWR VPWR genblk1_o3_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_533_ clknet_3_2_0_clk _026_ _045_ VGND VGND VPWR VPWR genblk1_o5_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_534_ clknet_3_2_0_clk genblk1_o5_c_dcsa_dhsum2 _046_ VGND VGND VPWR VPWR genblk1_o4_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_535_ clknet_3_2_0_clk _027_ _047_ VGND VGND VPWR VPWR genblk1_o6_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_536_ clknet_3_2_0_clk genblk1_o6_c_dcsa_dhsum2 _048_ VGND VGND VPWR VPWR genblk1_o5_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_537_ clknet_3_2_0_clk _028_ _049_ VGND VGND VPWR VPWR genblk1_o7_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_538_ clknet_3_2_0_clk genblk1_o7_c_dcsa_dhsum2 _050_ VGND VGND VPWR VPWR genblk1_o6_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_539_ clknet_3_3_0_clk _029_ _051_ VGND VGND VPWR VPWR genblk1_o8_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_540_ clknet_3_2_0_clk genblk1_o8_c_dcsa_dhsum2 _052_ VGND VGND VPWR VPWR genblk1_o7_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_541_ clknet_3_3_0_clk _030_ _053_ VGND VGND VPWR VPWR genblk1_o9_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_542_ clknet_3_3_0_clk genblk1_o9_c_dcsa_dhsum2 _054_ VGND VGND VPWR VPWR genblk1_o8_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_543_ clknet_3_6_0_clk _001_ _055_ VGND VGND VPWR VPWR genblk1_o10_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_544_ clknet_3_3_0_clk genblk1_o10_c_dcsa_dhsum2 _056_ VGND VGND VPWR VPWR genblk1_o10_c_dcsa_dsum
+ sky130_fd_sc_hd__dfrtp_1
X_545_ clknet_3_6_0_clk _002_ _057_ VGND VGND VPWR VPWR genblk1_o11_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_546_ clknet_3_3_0_clk genblk1_o11_c_dcsa_dhsum2 _058_ VGND VGND VPWR VPWR genblk1_o10_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_547_ clknet_3_3_0_clk _003_ _059_ VGND VGND VPWR VPWR genblk1_o12_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_548_ clknet_3_2_0_clk genblk1_o12_c_dcsa_dhsum2 _060_ VGND VGND VPWR VPWR genblk1_o11_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_549_ clknet_3_1_0_clk _004_ _061_ VGND VGND VPWR VPWR genblk1_o13_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_550_ clknet_3_1_0_clk genblk1_o13_c_dcsa_dhsum2 _062_ VGND VGND VPWR VPWR genblk1_o12_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_551_ clknet_3_1_0_clk _005_ _063_ VGND VGND VPWR VPWR genblk1_o14_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_552_ clknet_3_1_0_clk genblk1_o14_c_dcsa_dhsum2 _064_ VGND VGND VPWR VPWR genblk1_o13_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_553_ clknet_3_4_0_clk _006_ _065_ VGND VGND VPWR VPWR genblk1_o15_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_554_ clknet_3_4_0_clk genblk1_o15_c_dcsa_dhsum2 _066_ VGND VGND VPWR VPWR genblk1_o14_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_555_ clknet_3_4_0_clk _007_ _067_ VGND VGND VPWR VPWR genblk1_o16_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_556_ clknet_3_4_0_clk genblk1_o16_c_dcsa_dhsum2 _068_ VGND VGND VPWR VPWR genblk1_o15_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_557_ clknet_3_5_0_clk _008_ _069_ VGND VGND VPWR VPWR genblk1_o17_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_558_ clknet_3_4_0_clk genblk1_o17_c_dcsa_dhsum2 _070_ VGND VGND VPWR VPWR genblk1_o16_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_559_ clknet_3_6_0_clk _009_ _071_ VGND VGND VPWR VPWR genblk1_o18_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_560_ clknet_3_6_0_clk genblk1_o18_c_dcsa_dhsum2 _072_ VGND VGND VPWR VPWR genblk1_o17_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_561_ clknet_3_7_0_clk _010_ _073_ VGND VGND VPWR VPWR genblk1_o19_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_562_ clknet_3_6_0_clk genblk1_o19_c_dcsa_dhsum2 _074_ VGND VGND VPWR VPWR genblk1_o18_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_563_ clknet_3_6_0_clk _012_ _075_ VGND VGND VPWR VPWR genblk1_o20_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_564_ clknet_3_6_0_clk genblk1_o20_c_dcsa_dhsum2 _076_ VGND VGND VPWR VPWR genblk1_o19_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_565_ clknet_3_6_0_clk _013_ _077_ VGND VGND VPWR VPWR genblk1_o21_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_566_ clknet_3_7_0_clk genblk1_o21_c_dcsa_dhsum2 _078_ VGND VGND VPWR VPWR genblk1_o20_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_567_ clknet_3_7_0_clk _014_ _079_ VGND VGND VPWR VPWR genblk1_o22_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_568_ clknet_3_7_0_clk genblk1_o22_c_dcsa_dhsum2 _080_ VGND VGND VPWR VPWR genblk1_o21_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_569_ clknet_3_7_0_clk _015_ _081_ VGND VGND VPWR VPWR genblk1_o23_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_570_ clknet_3_7_0_clk genblk1_o23_c_dcsa_dhsum2 _082_ VGND VGND VPWR VPWR genblk1_o22_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_571_ clknet_3_7_0_clk _016_ _083_ VGND VGND VPWR VPWR genblk1_o24_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_572_ clknet_3_7_0_clk genblk1_o24_c_dcsa_dhsum2 _084_ VGND VGND VPWR VPWR genblk1_o23_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_573_ clknet_3_5_0_clk _017_ _085_ VGND VGND VPWR VPWR genblk1_o25_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_574_ clknet_3_7_0_clk genblk1_o25_c_dcsa_dhsum2 _086_ VGND VGND VPWR VPWR genblk1_o24_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_575_ clknet_3_5_0_clk _018_ _087_ VGND VGND VPWR VPWR genblk1_o26_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_576_ clknet_3_5_0_clk genblk1_o26_c_dcsa_dhsum2 _088_ VGND VGND VPWR VPWR genblk1_o25_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_577_ clknet_3_5_0_clk _019_ _089_ VGND VGND VPWR VPWR genblk1_o27_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_578_ clknet_3_5_0_clk genblk1_o27_c_dcsa_dhsum2 _090_ VGND VGND VPWR VPWR genblk1_o26_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_579_ clknet_3_5_0_clk _020_ _091_ VGND VGND VPWR VPWR genblk1_o28_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_580_ clknet_3_5_0_clk genblk1_o28_c_dcsa_dhsum2 _092_ VGND VGND VPWR VPWR genblk1_o27_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_581_ clknet_3_5_0_clk _021_ _093_ VGND VGND VPWR VPWR genblk1_o29_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_582_ clknet_3_5_0_clk genblk1_o29_c_dcsa_dhsum2 _094_ VGND VGND VPWR VPWR genblk1_o28_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
X_583_ clknet_3_4_0_clk _023_ _095_ VGND VGND VPWR VPWR genblk1_o30_c_dcsa_dsc
+ sky130_fd_sc_hd__dfrtp_1
X_584_ clknet_3_4_0_clk genblk1_o30_c_dcsa_dhsum2 _096_ VGND VGND VPWR VPWR genblk1_o29_c_dcsa_dy
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_0_0_clk clknet_1_0_0_clk VGND VGND VPWR VPWR clknet_2_0_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_clk clknet_1_0_0_clk VGND VGND VPWR VPWR clknet_2_1_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_2_0_clk clknet_1_1_0_clk VGND VGND VPWR VPWR clknet_2_2_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_3_0_clk clknet_1_1_0_clk VGND VGND VPWR VPWR clknet_2_3_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_0_0_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_1_0_clk clknet_2_0_0_clk VGND VGND VPWR VPWR clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_2_0_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_3_0_clk clknet_2_1_0_clk VGND VGND VPWR VPWR clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_4_0_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_5_0_clk clknet_2_2_0_clk VGND VGND VPWR VPWR clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_6_0_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_7_0_clk clknet_2_3_0_clk VGND VGND VPWR VPWR clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_2
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
Xinput10 x[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput11 x[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput12 x[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput13 x[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput14 x[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput15 x[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput16 x[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput17 x[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput18 x[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput19 x[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xinput2 x[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xinput20 x[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput21 x[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput22 x[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput23 x[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput24 x[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput25 x[30] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 x[31] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput27 x[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput28 x[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput29 x[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
Xinput3 x[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
Xinput30 x[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput31 x[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput32 x[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput33 x[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput34 y VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput4 x[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xinput5 x[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
Xinput6 x[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
Xinput7 x[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
Xinput8 x[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
Xinput9 x[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xoutput35 net35 VGND VGND VPWR VPWR p sky130_fd_sc_hd__buf_2
**.ends
.end
